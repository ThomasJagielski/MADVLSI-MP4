magic
tech sky130A
magscale 1 2
timestamp 1617356490
<< error_p >>
rect 5953 0 6000 3200
rect 6600 0 7200 3200
rect 7800 0 8400 3200
rect 9000 0 9600 3200
rect 10200 0 10800 3200
rect 11400 0 12000 3200
rect 12600 0 13200 3200
rect 13800 0 14400 3200
rect 15000 0 15600 3200
rect 16200 0 16800 3200
rect 17400 0 18000 3200
rect 18600 0 19200 3200
rect 19800 0 19847 3200
rect 5953 -4000 6000 -800
rect 6600 -4000 7200 -800
rect 7800 -4000 8400 -800
rect 9000 -4000 9600 -800
rect 10200 -4000 10800 -800
rect 11400 -4000 12000 -800
rect 12600 -4000 13200 -800
rect 13800 -4000 14400 -800
rect 15000 -4000 15600 -800
rect 16200 -4000 16800 -800
rect 17400 -4000 18000 -800
rect 18600 -4000 19200 -800
rect 19800 -4000 19847 -800
rect 5953 -8000 6000 -4800
rect 6600 -8000 7200 -4800
rect 7800 -8000 8400 -4800
rect 9000 -8000 9600 -4800
rect 10200 -8000 10800 -4800
rect 11400 -8000 12000 -4800
rect 12600 -8000 13200 -4800
rect 13800 -8000 14400 -4800
rect 15000 -8000 15600 -4800
rect 16200 -8000 16800 -4800
rect 17400 -8000 18000 -4800
rect 18600 -8000 19200 -4800
rect 19800 -8000 19847 -4800
<< nmos >>
rect -2400 0 -1800 3200
rect -1200 0 -600 3200
rect 0 0 600 3200
rect 1200 0 1800 3200
rect 4800 0 5400 3200
rect 6000 0 6600 3200
rect 7200 0 7800 3200
rect 8400 0 9000 3200
rect 9600 0 10200 3200
rect 10800 0 11400 3200
rect 12000 0 12600 3200
rect 13200 0 13800 3200
rect 14400 0 15000 3200
rect 15600 0 16200 3200
rect 16800 0 17400 3200
rect 18000 0 18600 3200
rect 19200 0 19800 3200
rect 20400 0 21000 3200
rect 21600 0 22200 3200
rect -2400 -4000 -1800 -800
rect -1200 -4000 -600 -800
rect 0 -4000 600 -800
rect 1200 -4000 1800 -800
rect 4800 -4000 5400 -800
rect 6000 -4000 6600 -800
rect 7200 -4000 7800 -800
rect 8400 -4000 9000 -800
rect 9600 -4000 10200 -800
rect 10800 -4000 11400 -800
rect 12000 -4000 12600 -800
rect 13200 -4000 13800 -800
rect 14400 -4000 15000 -800
rect 15600 -4000 16200 -800
rect 16800 -4000 17400 -800
rect 18000 -4000 18600 -800
rect 19200 -4000 19800 -800
rect 20400 -4000 21000 -800
rect 21600 -4000 22200 -800
rect -2400 -8000 -1800 -4800
rect -1200 -8000 -600 -4800
rect 0 -8000 600 -4800
rect 1200 -8000 1800 -4800
rect 4800 -8000 5400 -4800
rect 6000 -8000 6600 -4800
rect 7200 -8000 7800 -4800
rect 8400 -8000 9000 -4800
rect 9600 -8000 10200 -4800
rect 10800 -8000 11400 -4800
rect 12000 -8000 12600 -4800
rect 13200 -8000 13800 -4800
rect 14400 -8000 15000 -4800
rect 15600 -8000 16200 -4800
rect 16800 -8000 17400 -4800
rect 18000 -8000 18600 -4800
rect 19200 -8000 19800 -4800
rect 20400 -8000 21000 -4800
rect 21600 -8000 22200 -4800
<< ndiff >>
rect -3000 3170 -2400 3200
rect -3000 30 -2970 3170
rect -2430 30 -2400 3170
rect -3000 0 -2400 30
rect -1800 3170 -1200 3200
rect -1800 30 -1770 3170
rect -1230 30 -1200 3170
rect -1800 0 -1200 30
rect -600 3170 0 3200
rect -600 30 -570 3170
rect -30 30 0 3170
rect -600 0 0 30
rect 600 3170 1200 3200
rect 600 30 630 3170
rect 1170 30 1200 3170
rect 600 0 1200 30
rect 1800 3170 2400 3200
rect 1800 30 1830 3170
rect 2370 30 2400 3170
rect 1800 0 2400 30
rect 3000 0 4800 3200
rect 5400 3170 6000 3200
rect 5400 30 5430 3170
rect 5970 30 6000 3170
rect 5400 0 6000 30
rect 6600 3170 7200 3200
rect 6600 30 6630 3170
rect 7170 30 7200 3170
rect 6600 0 7200 30
rect 7800 3170 8400 3200
rect 7800 30 7830 3170
rect 8370 30 8400 3170
rect 7800 0 8400 30
rect 9000 3170 9600 3200
rect 9000 30 9030 3170
rect 9570 30 9600 3170
rect 9000 0 9600 30
rect 10200 3170 10800 3200
rect 10200 30 10230 3170
rect 10770 30 10800 3170
rect 10200 0 10800 30
rect 11400 3170 12000 3200
rect 11400 30 11430 3170
rect 11970 30 12000 3170
rect 11400 0 12000 30
rect 12600 3170 13200 3200
rect 12600 30 12630 3170
rect 13170 30 13200 3170
rect 12600 0 13200 30
rect 13800 3170 14400 3200
rect 13800 30 13830 3170
rect 14370 30 14400 3170
rect 13800 0 14400 30
rect 15000 3170 15600 3200
rect 15000 30 15030 3170
rect 15570 30 15600 3170
rect 15000 0 15600 30
rect 16200 3170 16800 3200
rect 16200 30 16230 3170
rect 16770 30 16800 3170
rect 16200 0 16800 30
rect 17400 3170 18000 3200
rect 17400 30 17430 3170
rect 17970 30 18000 3170
rect 17400 0 18000 30
rect 18600 3170 19200 3200
rect 18600 30 18630 3170
rect 19170 30 19200 3170
rect 18600 0 19200 30
rect 19800 3170 20400 3200
rect 19800 30 19830 3170
rect 20370 30 20400 3170
rect 19800 0 20400 30
rect 21000 3170 21600 3200
rect 21000 30 21030 3170
rect 21570 30 21600 3170
rect 21000 0 21600 30
rect 22200 3170 22800 3200
rect 22200 30 22230 3170
rect 22770 30 22800 3170
rect 22200 0 22800 30
rect -3000 -830 -2400 -800
rect -3000 -3970 -2970 -830
rect -2430 -3970 -2400 -830
rect -3000 -4000 -2400 -3970
rect -1800 -830 -1200 -800
rect -1800 -3970 -1770 -830
rect -1230 -3970 -1200 -830
rect -1800 -4000 -1200 -3970
rect -600 -830 0 -800
rect -600 -3970 -570 -830
rect -30 -3970 0 -830
rect -600 -4000 0 -3970
rect 600 -830 1200 -800
rect 600 -3970 630 -830
rect 1170 -3970 1200 -830
rect 600 -4000 1200 -3970
rect 1800 -830 2400 -800
rect 1800 -3970 1830 -830
rect 2370 -3970 2400 -830
rect 1800 -4000 2400 -3970
rect 3000 -4000 4800 -800
rect 5400 -830 6000 -800
rect 5400 -3970 5430 -830
rect 5970 -3970 6000 -830
rect 5400 -4000 6000 -3970
rect 6600 -830 7200 -800
rect 6600 -3970 6630 -830
rect 7170 -3970 7200 -830
rect 6600 -4000 7200 -3970
rect 7800 -830 8400 -800
rect 7800 -3970 7830 -830
rect 8370 -3970 8400 -830
rect 7800 -4000 8400 -3970
rect 9000 -830 9600 -800
rect 9000 -3970 9030 -830
rect 9570 -3970 9600 -830
rect 9000 -4000 9600 -3970
rect 10200 -830 10800 -800
rect 10200 -3970 10230 -830
rect 10770 -3970 10800 -830
rect 10200 -4000 10800 -3970
rect 11400 -830 12000 -800
rect 11400 -3970 11430 -830
rect 11970 -3970 12000 -830
rect 11400 -4000 12000 -3970
rect 12600 -830 13200 -800
rect 12600 -3970 12630 -830
rect 13170 -3970 13200 -830
rect 12600 -4000 13200 -3970
rect 13800 -830 14400 -800
rect 13800 -3970 13830 -830
rect 14370 -3970 14400 -830
rect 13800 -4000 14400 -3970
rect 15000 -830 15600 -800
rect 15000 -3970 15030 -830
rect 15570 -3970 15600 -830
rect 15000 -4000 15600 -3970
rect 16200 -830 16800 -800
rect 16200 -3970 16230 -830
rect 16770 -3970 16800 -830
rect 16200 -4000 16800 -3970
rect 17400 -830 18000 -800
rect 17400 -3970 17430 -830
rect 17970 -3970 18000 -830
rect 17400 -4000 18000 -3970
rect 18600 -830 19200 -800
rect 18600 -3970 18630 -830
rect 19170 -3970 19200 -830
rect 18600 -4000 19200 -3970
rect 19800 -830 20400 -800
rect 19800 -3970 19830 -830
rect 20370 -3970 20400 -830
rect 19800 -4000 20400 -3970
rect 21000 -830 21600 -800
rect 21000 -3970 21030 -830
rect 21570 -3970 21600 -830
rect 21000 -4000 21600 -3970
rect 22200 -830 22800 -800
rect 22200 -3970 22230 -830
rect 22770 -3970 22800 -830
rect 22200 -4000 22800 -3970
rect -3000 -4830 -2400 -4800
rect -3000 -7970 -2970 -4830
rect -2430 -7970 -2400 -4830
rect -3000 -8000 -2400 -7970
rect -1800 -4830 -1200 -4800
rect -1800 -7970 -1770 -4830
rect -1230 -7970 -1200 -4830
rect -1800 -8000 -1200 -7970
rect -600 -4830 0 -4800
rect -600 -7970 -570 -4830
rect -30 -7970 0 -4830
rect -600 -8000 0 -7970
rect 600 -4830 1200 -4800
rect 600 -7970 630 -4830
rect 1170 -7970 1200 -4830
rect 600 -8000 1200 -7970
rect 1800 -4830 2400 -4800
rect 1800 -7970 1830 -4830
rect 2370 -7970 2400 -4830
rect 1800 -8000 2400 -7970
rect 3000 -8000 4800 -4800
rect 5400 -4830 6000 -4800
rect 5400 -7970 5430 -4830
rect 5970 -7970 6000 -4830
rect 5400 -8000 6000 -7970
rect 6600 -4830 7200 -4800
rect 6600 -7970 6630 -4830
rect 7170 -7970 7200 -4830
rect 6600 -8000 7200 -7970
rect 7800 -4830 8400 -4800
rect 7800 -7970 7830 -4830
rect 8370 -7970 8400 -4830
rect 7800 -8000 8400 -7970
rect 9000 -4830 9600 -4800
rect 9000 -7970 9030 -4830
rect 9570 -7970 9600 -4830
rect 9000 -8000 9600 -7970
rect 10200 -4830 10800 -4800
rect 10200 -7970 10230 -4830
rect 10770 -7970 10800 -4830
rect 10200 -8000 10800 -7970
rect 11400 -4830 12000 -4800
rect 11400 -7970 11430 -4830
rect 11970 -7970 12000 -4830
rect 11400 -8000 12000 -7970
rect 12600 -4830 13200 -4800
rect 12600 -7970 12630 -4830
rect 13170 -7970 13200 -4830
rect 12600 -8000 13200 -7970
rect 13800 -4830 14400 -4800
rect 13800 -7970 13830 -4830
rect 14370 -7970 14400 -4830
rect 13800 -8000 14400 -7970
rect 15000 -4830 15600 -4800
rect 15000 -7970 15030 -4830
rect 15570 -7970 15600 -4830
rect 15000 -8000 15600 -7970
rect 16200 -4830 16800 -4800
rect 16200 -7970 16230 -4830
rect 16770 -7970 16800 -4830
rect 16200 -8000 16800 -7970
rect 17400 -4830 18000 -4800
rect 17400 -7970 17430 -4830
rect 17970 -7970 18000 -4830
rect 17400 -8000 18000 -7970
rect 18600 -4830 19200 -4800
rect 18600 -7970 18630 -4830
rect 19170 -7970 19200 -4830
rect 18600 -8000 19200 -7970
rect 19800 -4830 20400 -4800
rect 19800 -7970 19830 -4830
rect 20370 -7970 20400 -4830
rect 19800 -8000 20400 -7970
rect 21000 -4830 21600 -4800
rect 21000 -7970 21030 -4830
rect 21570 -7970 21600 -4830
rect 21000 -8000 21600 -7970
rect 22200 -4830 22800 -4800
rect 22200 -7970 22230 -4830
rect 22770 -7970 22800 -4830
rect 22200 -8000 22800 -7970
<< ndiffc >>
rect -2970 30 -2430 3170
rect -1770 30 -1230 3170
rect -570 30 -30 3170
rect 630 30 1170 3170
rect 1830 30 2370 3170
rect 5430 30 5970 3170
rect 6630 30 7170 3170
rect 7830 30 8370 3170
rect 9030 30 9570 3170
rect 10230 30 10770 3170
rect 11430 30 11970 3170
rect 12630 30 13170 3170
rect 13830 30 14370 3170
rect 15030 30 15570 3170
rect 16230 30 16770 3170
rect 17430 30 17970 3170
rect 18630 30 19170 3170
rect 19830 30 20370 3170
rect 21030 30 21570 3170
rect 22230 30 22770 3170
rect -2970 -3970 -2430 -830
rect -1770 -3970 -1230 -830
rect -570 -3970 -30 -830
rect 630 -3970 1170 -830
rect 1830 -3970 2370 -830
rect 5430 -3970 5970 -830
rect 6630 -3970 7170 -830
rect 7830 -3970 8370 -830
rect 9030 -3970 9570 -830
rect 10230 -3970 10770 -830
rect 11430 -3970 11970 -830
rect 12630 -3970 13170 -830
rect 13830 -3970 14370 -830
rect 15030 -3970 15570 -830
rect 16230 -3970 16770 -830
rect 17430 -3970 17970 -830
rect 18630 -3970 19170 -830
rect 19830 -3970 20370 -830
rect 21030 -3970 21570 -830
rect 22230 -3970 22770 -830
rect -2970 -7970 -2430 -4830
rect -1770 -7970 -1230 -4830
rect -570 -7970 -30 -4830
rect 630 -7970 1170 -4830
rect 1830 -7970 2370 -4830
rect 5430 -7970 5970 -4830
rect 6630 -7970 7170 -4830
rect 7830 -7970 8370 -4830
rect 9030 -7970 9570 -4830
rect 10230 -7970 10770 -4830
rect 11430 -7970 11970 -4830
rect 12630 -7970 13170 -4830
rect 13830 -7970 14370 -4830
rect 15030 -7970 15570 -4830
rect 16230 -7970 16770 -4830
rect 17430 -7970 17970 -4830
rect 18630 -7970 19170 -4830
rect 19830 -7970 20370 -4830
rect 21030 -7970 21570 -4830
rect 22230 -7970 22770 -4830
<< psubdiff >>
rect -3600 3170 -3000 3200
rect -3600 30 -3570 3170
rect -3030 30 -3000 3170
rect -3600 0 -3000 30
rect 2400 3170 3000 3200
rect 2400 30 2430 3170
rect 2970 30 3000 3170
rect 2400 0 3000 30
rect 22800 3170 23400 3200
rect 22800 30 22830 3170
rect 23370 30 23400 3170
rect 22800 0 23400 30
rect -3600 -830 -3000 -800
rect -3600 -3970 -3570 -830
rect -3030 -3970 -3000 -830
rect -3600 -4000 -3000 -3970
rect 2400 -830 3000 -800
rect 2400 -3970 2430 -830
rect 2970 -3970 3000 -830
rect 2400 -4000 3000 -3970
rect 22800 -830 23400 -800
rect 22800 -3970 22830 -830
rect 23370 -3970 23400 -830
rect 22800 -4000 23400 -3970
rect -3600 -4830 -3000 -4800
rect -3600 -7970 -3570 -4830
rect -3030 -7970 -3000 -4830
rect -3600 -8000 -3000 -7970
rect 2400 -4830 3000 -4800
rect 2400 -7970 2430 -4830
rect 2970 -7970 3000 -4830
rect 2400 -8000 3000 -7970
rect 22800 -4830 23400 -4800
rect 22800 -7970 22830 -4830
rect 23370 -7970 23400 -4830
rect 22800 -8000 23400 -7970
<< psubdiffcont >>
rect -3570 30 -3030 3170
rect 2430 30 2970 3170
rect 22830 30 23370 3170
rect -3570 -3970 -3030 -830
rect 2430 -3970 2970 -830
rect 22830 -3970 23370 -830
rect -3570 -7970 -3030 -4830
rect 2430 -7970 2970 -4830
rect 22830 -7970 23370 -4830
<< poly >>
rect 19720 3370 19800 3390
rect 19720 3330 19740 3370
rect 19780 3330 19800 3370
rect 19720 3310 19800 3330
rect -2740 3290 -2660 3310
rect -2740 3260 -2720 3290
rect -2990 3250 -2720 3260
rect -2680 3260 -2660 3290
rect -1540 3290 -1460 3310
rect -1540 3260 -1520 3290
rect -2680 3250 -1520 3260
rect -1480 3260 -1460 3290
rect 0 3280 19800 3310
rect -1480 3250 -600 3260
rect -2990 3230 -600 3250
rect -2400 3200 -1800 3230
rect -1200 3200 -600 3230
rect 0 3200 600 3280
rect 1200 3200 1800 3280
rect 4800 3200 5400 3230
rect 6000 3200 6600 3280
rect 7200 3200 7800 3230
rect 8400 3200 9000 3280
rect 9600 3200 10200 3230
rect 10800 3200 11400 3280
rect 12000 3200 12600 3230
rect 13200 3200 13800 3280
rect 14400 3200 15000 3230
rect 15600 3200 16200 3280
rect 16800 3200 17400 3230
rect 18000 3200 18600 3280
rect 19200 3200 19800 3280
rect 21240 3290 21320 3310
rect 21240 3260 21260 3290
rect 20400 3250 21260 3260
rect 21300 3260 21320 3290
rect 22460 3290 22540 3310
rect 22460 3260 22480 3290
rect 21300 3250 22480 3260
rect 22520 3260 22540 3290
rect 22520 3250 22790 3260
rect 20400 3230 22790 3250
rect 20400 3200 21000 3230
rect 21600 3200 22200 3230
rect -2400 -30 -1800 0
rect -1200 -30 -600 0
rect 0 -30 600 0
rect 1200 -30 1800 0
rect 4800 -30 5400 0
rect 6000 -30 6600 0
rect 7200 -30 7800 0
rect 8400 -30 9000 0
rect 9600 -30 10200 0
rect 10800 -30 11400 0
rect 12000 -30 12600 0
rect 13200 -30 13800 0
rect 14400 -30 15000 0
rect 15600 -30 16200 0
rect 16800 -30 17400 0
rect 18000 -30 18600 0
rect 19200 -30 19800 0
rect 20400 -30 21000 0
rect 21600 -30 22200 0
rect 5060 -50 5140 -30
rect 5060 -90 5080 -50
rect 5120 -90 5140 -50
rect 5060 -110 5140 -90
rect 7460 -50 7540 -30
rect 7460 -90 7480 -50
rect 7520 -90 7540 -50
rect 7460 -110 7540 -90
rect 9860 -50 9940 -30
rect 9860 -90 9880 -50
rect 9920 -90 9940 -50
rect 9860 -110 9940 -90
rect 12260 -50 12340 -30
rect 12260 -90 12280 -50
rect 12320 -90 12340 -50
rect 12260 -110 12340 -90
rect 14660 -50 14740 -30
rect 14660 -90 14680 -50
rect 14720 -90 14740 -50
rect 14660 -110 14740 -90
rect 17060 -50 17140 -30
rect 17060 -90 17080 -50
rect 17120 -90 17140 -50
rect 17060 -110 17140 -90
rect 7200 -560 7800 -530
rect 7200 -660 7230 -560
rect 0 -690 7230 -660
rect 7770 -660 7800 -560
rect 13200 -560 13800 -530
rect 13200 -660 13230 -560
rect 7770 -690 13230 -660
rect 13770 -660 13800 -560
rect 18300 -660 18330 -30
rect 13770 -690 18600 -660
rect -2740 -710 -2660 -690
rect -2740 -740 -2720 -710
rect -2990 -750 -2720 -740
rect -2680 -740 -2660 -710
rect -1540 -710 -1460 -690
rect -1540 -740 -1520 -710
rect -2680 -750 -1520 -740
rect -1480 -740 -1460 -710
rect -1480 -750 -600 -740
rect -2990 -770 -600 -750
rect -2400 -800 -1800 -770
rect -1200 -800 -600 -770
rect 0 -800 600 -690
rect 1200 -800 1800 -690
rect 4800 -800 5400 -690
rect 6000 -800 6600 -690
rect 7460 -710 7540 -690
rect 7460 -750 7480 -710
rect 7520 -750 7540 -710
rect 7460 -770 7540 -750
rect 7200 -800 7800 -770
rect 8400 -800 9000 -690
rect 9600 -800 10200 -690
rect 10800 -800 11400 -690
rect 12000 -800 12600 -690
rect 13460 -710 13540 -690
rect 13460 -750 13480 -710
rect 13520 -750 13540 -710
rect 13460 -770 13540 -750
rect 13200 -800 13800 -770
rect 14400 -800 15000 -690
rect 15600 -800 16200 -690
rect 16800 -800 17400 -690
rect 18000 -800 18600 -690
rect 20060 -710 20140 -690
rect 20060 -740 20080 -710
rect 19200 -750 20080 -740
rect 20120 -740 20140 -710
rect 21260 -710 21340 -690
rect 21260 -740 21280 -710
rect 20120 -750 21280 -740
rect 21320 -740 21340 -710
rect 22460 -710 22540 -690
rect 22460 -740 22480 -710
rect 21320 -750 22480 -740
rect 22520 -740 22540 -710
rect 22520 -750 22790 -740
rect 19200 -770 22790 -750
rect 19200 -800 19800 -770
rect 20400 -800 21000 -770
rect 21600 -800 22200 -770
rect -2400 -4030 -1800 -4000
rect -1200 -4030 -600 -4000
rect 0 -4030 600 -4000
rect 1200 -4030 1800 -4000
rect 4800 -4030 5400 -4000
rect 6000 -4030 6600 -4000
rect 7200 -4030 7800 -4000
rect 8400 -4030 9000 -4000
rect 9600 -4030 10200 -4000
rect 10800 -4030 11400 -4000
rect 12000 -4030 12600 -4000
rect 13200 -4030 13800 -4000
rect 14400 -4030 15000 -4000
rect 15600 -4030 16200 -4000
rect 16800 -4030 17400 -4000
rect 18000 -4030 18600 -4000
rect 19200 -4030 19800 -4000
rect 20400 -4030 21000 -4000
rect 21600 -4030 22200 -4000
rect 1070 -4050 1150 -4030
rect 1070 -4090 1090 -4050
rect 1130 -4090 1150 -4050
rect 1070 -4110 1150 -4090
rect 9260 -4050 9340 -4030
rect 9260 -4090 9280 -4050
rect 9320 -4090 9340 -4050
rect 9260 -4110 9340 -4090
rect 15050 -4050 15130 -4030
rect 15050 -4090 15070 -4050
rect 15110 -4090 15130 -4050
rect 15050 -4110 15130 -4090
rect 17450 -4050 17530 -4030
rect 17450 -4090 17470 -4050
rect 17510 -4090 17530 -4050
rect 17450 -4110 17530 -4090
rect 1070 -4670 1100 -4110
rect 1070 -4690 1150 -4670
rect 1070 -4730 1090 -4690
rect 1130 -4730 1150 -4690
rect 1070 -4750 1150 -4730
rect 9260 -4690 9290 -4110
rect 15050 -4590 15080 -4110
rect 15050 -4610 15130 -4590
rect 15050 -4650 15070 -4610
rect 15110 -4650 15130 -4610
rect 15050 -4670 15130 -4650
rect 17450 -4680 17480 -4110
rect 9260 -4710 9340 -4690
rect 9260 -4750 9280 -4710
rect 9320 -4750 9340 -4710
rect 9260 -4770 9340 -4750
rect 17450 -4700 17530 -4680
rect 17450 -4740 17470 -4700
rect 17510 -4740 17530 -4700
rect 17450 -4760 17530 -4740
rect -2400 -4800 -1800 -4770
rect -1200 -4800 -600 -4770
rect 0 -4800 600 -4770
rect 1200 -4800 1800 -4770
rect 4800 -4800 5400 -4770
rect 6000 -4800 6600 -4770
rect 7200 -4800 7800 -4770
rect 8400 -4800 9000 -4770
rect 9600 -4800 10200 -4770
rect 10800 -4800 11400 -4770
rect 12000 -4800 12600 -4770
rect 13200 -4800 13800 -4770
rect 14400 -4800 15000 -4770
rect 15600 -4800 16200 -4770
rect 16800 -4800 17400 -4770
rect 18000 -4800 18600 -4770
rect 19200 -4800 19800 -4770
rect 20400 -4800 21000 -4770
rect 21600 -4800 22200 -4770
rect -2400 -8030 -1800 -8000
rect -1200 -8030 -600 -8000
rect 0 -8030 600 -8000
rect 1200 -8030 1800 -8000
rect 4800 -8030 5400 -8000
rect 6000 -8030 6600 -8000
rect 7200 -8030 7800 -8000
rect 8400 -8030 9000 -8000
rect 9600 -8030 10200 -8000
rect 10800 -8030 11400 -8000
rect 12000 -8030 12600 -8000
rect 13200 -8030 13800 -8000
rect 14400 -8030 15000 -8000
rect 15600 -8030 16200 -8000
rect 16800 -8030 17400 -8000
rect 18000 -8030 18600 -8000
rect 19200 -8030 19800 -8000
rect 20400 -8030 21000 -8000
rect 21600 -8030 22200 -8000
rect -2990 -8050 1800 -8030
rect -2990 -8060 -2720 -8050
rect -2740 -8090 -2720 -8060
rect -2680 -8060 -1520 -8050
rect -2680 -8090 -2660 -8060
rect -2740 -8110 -2660 -8090
rect -1540 -8090 -1520 -8060
rect -1480 -8060 -320 -8050
rect -1480 -8090 -1460 -8060
rect -1540 -8110 -1460 -8090
rect -340 -8090 -320 -8060
rect -280 -8060 880 -8050
rect -280 -8090 -260 -8060
rect -340 -8110 -260 -8090
rect 860 -8090 880 -8060
rect 920 -8060 1800 -8050
rect 6260 -8050 6340 -8030
rect 920 -8090 940 -8060
rect 860 -8110 940 -8090
rect 6260 -8090 6280 -8050
rect 6320 -8090 6340 -8050
rect 6260 -8110 6340 -8090
rect 7460 -8050 7540 -8030
rect 7460 -8090 7480 -8050
rect 7520 -8090 7540 -8050
rect 7460 -8110 7540 -8090
rect 8660 -8050 8740 -8030
rect 8660 -8090 8680 -8050
rect 8720 -8090 8740 -8050
rect 8660 -8110 8740 -8090
rect 9860 -8050 9940 -8030
rect 9860 -8090 9880 -8050
rect 9920 -8090 9940 -8050
rect 9860 -8110 9940 -8090
rect 11060 -8050 11140 -8030
rect 11060 -8090 11080 -8050
rect 11120 -8090 11140 -8050
rect 11060 -8110 11140 -8090
rect 12260 -8050 12340 -8030
rect 12260 -8090 12280 -8050
rect 12320 -8090 12340 -8050
rect 12260 -8110 12340 -8090
rect 13460 -8050 13540 -8030
rect 13460 -8090 13480 -8050
rect 13520 -8090 13540 -8050
rect 13460 -8110 13540 -8090
rect 14660 -8050 14740 -8030
rect 14660 -8090 14680 -8050
rect 14720 -8090 14740 -8050
rect 14660 -8110 14740 -8090
rect 15860 -8050 15940 -8030
rect 15860 -8090 15880 -8050
rect 15920 -8090 15940 -8050
rect 16800 -8050 22790 -8030
rect 16800 -8060 17680 -8050
rect 15860 -8110 15940 -8090
rect 17660 -8090 17680 -8060
rect 17720 -8060 18880 -8050
rect 17720 -8090 17740 -8060
rect 17660 -8110 17740 -8090
rect 18860 -8090 18880 -8060
rect 18920 -8060 20080 -8050
rect 18920 -8090 18940 -8060
rect 18860 -8110 18940 -8090
rect 20060 -8090 20080 -8060
rect 20120 -8060 21280 -8050
rect 20120 -8090 20140 -8060
rect 20060 -8110 20140 -8090
rect 21260 -8090 21280 -8060
rect 21320 -8060 22480 -8050
rect 21320 -8090 21340 -8060
rect 21260 -8110 21340 -8090
rect 22460 -8090 22480 -8060
rect 22520 -8060 22790 -8050
rect 22520 -8090 22540 -8060
rect 22460 -8110 22540 -8090
<< polycont >>
rect 19740 3330 19780 3370
rect -2720 3250 -2680 3290
rect -1520 3250 -1480 3290
rect 21260 3250 21300 3290
rect 22480 3250 22520 3290
rect 5080 -90 5120 -50
rect 7480 -90 7520 -50
rect 9880 -90 9920 -50
rect 12280 -90 12320 -50
rect 14680 -90 14720 -50
rect 17080 -90 17120 -50
rect -2720 -750 -2680 -710
rect -1520 -750 -1480 -710
rect 7480 -750 7520 -710
rect 13480 -750 13520 -710
rect 20080 -750 20120 -710
rect 21280 -750 21320 -710
rect 22480 -750 22520 -710
rect 1090 -4090 1130 -4050
rect 9280 -4090 9320 -4050
rect 15070 -4090 15110 -4050
rect 17470 -4090 17510 -4050
rect 1090 -4730 1130 -4690
rect 15070 -4650 15110 -4610
rect 9280 -4750 9320 -4710
rect 17470 -4740 17510 -4700
rect -2720 -8090 -2680 -8050
rect -1520 -8090 -1480 -8050
rect -320 -8090 -280 -8050
rect 880 -8090 920 -8050
rect 6280 -8090 6320 -8050
rect 7480 -8090 7520 -8050
rect 8680 -8090 8720 -8050
rect 9880 -8090 9920 -8050
rect 11080 -8090 11120 -8050
rect 12280 -8090 12320 -8050
rect 13480 -8090 13520 -8050
rect 14680 -8090 14720 -8050
rect 15880 -8090 15920 -8050
rect 17680 -8090 17720 -8050
rect 18880 -8090 18920 -8050
rect 20080 -8090 20120 -8050
rect 21280 -8090 21320 -8050
rect 22480 -8090 22520 -8050
<< locali >>
rect 18610 3480 23400 3520
rect -2740 3290 -2660 3310
rect -2740 3250 -2720 3290
rect -2680 3250 -2660 3290
rect -2740 3230 -2660 3250
rect -1540 3290 -1460 3310
rect -1540 3250 -1520 3290
rect -1480 3250 -1460 3290
rect -1540 3230 -1460 3250
rect -2990 3190 -2410 3230
rect -3590 3170 -2410 3190
rect -3590 30 -3570 3170
rect -3030 30 -2970 3170
rect -2430 30 -2410 3170
rect -3590 10 -2410 30
rect -1790 3170 -1210 3230
rect -1790 30 -1770 3170
rect -1230 30 -1210 3170
rect -1790 10 -1210 30
rect -590 3170 -10 3190
rect -590 30 -570 3170
rect -30 30 -10 3170
rect -590 -40 -10 30
rect 610 3170 1190 3190
rect 610 30 630 3170
rect 1170 30 1190 3170
rect 610 10 1190 30
rect 1810 3170 2990 3190
rect 1810 30 1830 3170
rect 2370 30 2430 3170
rect 2970 30 2990 3170
rect 1810 10 2990 30
rect 5410 3170 5990 3190
rect 5410 30 5430 3170
rect 5970 30 5990 3170
rect 1810 -40 2390 10
rect -590 -80 2390 -40
rect 5060 -50 5140 -30
rect -2740 -710 -2660 -690
rect -2740 -750 -2720 -710
rect -2680 -750 -2660 -710
rect -2740 -770 -2660 -750
rect -1540 -710 -1460 -690
rect -1540 -750 -1520 -710
rect -1480 -750 -1460 -710
rect -1540 -770 -1460 -750
rect 880 -770 920 -80
rect 5060 -90 5080 -50
rect 5120 -90 5140 -50
rect 5410 -80 5990 30
rect 6610 3170 7190 3190
rect 6610 30 6630 3170
rect 7170 30 7190 3170
rect 6610 10 7190 30
rect 7810 3170 8390 3190
rect 7810 30 7830 3170
rect 8370 30 8390 3170
rect 7810 10 8390 30
rect 9010 3170 9590 3190
rect 9010 30 9030 3170
rect 9570 30 9590 3170
rect 7460 -50 7540 -30
rect 5060 -130 5140 -90
rect 5060 -170 5080 -130
rect 5120 -170 5140 -130
rect 5060 -190 5140 -170
rect 5680 -590 5720 -80
rect 7460 -90 7480 -50
rect 7520 -90 7540 -50
rect 9010 -80 9590 30
rect 10210 3170 10790 3190
rect 10210 30 10230 3170
rect 10770 30 10790 3170
rect 9860 -50 9940 -30
rect 7460 -130 7540 -90
rect 7460 -170 7480 -130
rect 7520 -170 7540 -130
rect 7460 -190 7540 -170
rect 1810 -630 5720 -590
rect 7200 -560 7800 -520
rect -2990 -810 -2410 -770
rect -3590 -830 -2410 -810
rect -3590 -3970 -3570 -830
rect -3030 -3970 -2970 -830
rect -2430 -3970 -2410 -830
rect -3590 -3990 -2410 -3970
rect -1790 -830 -1210 -770
rect -1790 -3970 -1770 -830
rect -1230 -3970 -1210 -830
rect -1790 -3990 -1210 -3970
rect -590 -830 -10 -810
rect -590 -3970 -570 -830
rect -30 -3970 -10 -830
rect -590 -4160 -10 -3970
rect 610 -830 1190 -770
rect 610 -3970 630 -830
rect 1170 -3970 1190 -830
rect 610 -4030 1190 -3970
rect 1810 -810 2390 -630
rect 7200 -680 7240 -560
rect 5410 -720 7240 -680
rect 7460 -630 7540 -610
rect 7460 -670 7480 -630
rect 7520 -670 7540 -630
rect 7460 -710 7540 -670
rect 1810 -830 2990 -810
rect 1810 -3970 1830 -830
rect 2370 -3970 2430 -830
rect 2970 -3970 2990 -830
rect 1810 -3990 2990 -3970
rect 5410 -830 5990 -720
rect 7460 -750 7480 -710
rect 7520 -750 7540 -710
rect 7760 -680 7800 -560
rect 9280 -680 9320 -80
rect 9860 -90 9880 -50
rect 9920 -90 9940 -50
rect 10210 -70 10790 30
rect 11410 3170 11990 3190
rect 11410 30 11430 3170
rect 11970 30 11990 3170
rect 11410 10 11990 30
rect 12610 3170 13190 3190
rect 12610 30 12630 3170
rect 13170 30 13190 3170
rect 12260 -50 12340 -30
rect 9860 -130 9940 -90
rect 9860 -170 9880 -130
rect 9920 -170 9940 -130
rect 9860 -190 9940 -170
rect 10480 -680 10520 -70
rect 12260 -90 12280 -50
rect 12320 -90 12340 -50
rect 12610 -70 13190 30
rect 13810 3170 14390 3190
rect 13810 30 13830 3170
rect 14370 30 14390 3170
rect 13810 10 14390 30
rect 15010 3170 15590 3190
rect 15010 30 15030 3170
rect 15570 30 15590 3170
rect 12260 -130 12340 -90
rect 12260 -170 12280 -130
rect 12320 -170 12340 -130
rect 12260 -190 12340 -170
rect 13150 -520 13190 -70
rect 14660 -50 14740 -30
rect 14660 -90 14680 -50
rect 14720 -90 14740 -50
rect 15010 -70 15590 30
rect 16210 3170 16790 3190
rect 16210 30 16230 3170
rect 16770 30 16790 3170
rect 16210 10 16790 30
rect 17410 3170 17990 3190
rect 17410 30 17430 3170
rect 17970 30 17990 3170
rect 17060 -50 17140 -30
rect 14660 -130 14740 -90
rect 14660 -170 14680 -130
rect 14720 -170 14740 -130
rect 14660 -190 14740 -170
rect 13150 -560 13800 -520
rect 13460 -630 13540 -610
rect 13460 -670 13480 -630
rect 13520 -670 13540 -630
rect 7760 -720 9590 -680
rect 7460 -770 7540 -750
rect 5410 -3970 5430 -830
rect 5970 -3970 5990 -830
rect 5410 -3990 5990 -3970
rect 6610 -830 7190 -810
rect 6610 -3970 6630 -830
rect 7170 -3970 7190 -830
rect 1070 -4050 1150 -4030
rect 1070 -4090 1090 -4050
rect 1130 -4090 1150 -4050
rect 1070 -4110 1150 -4090
rect 1810 -4160 2390 -3990
rect 6610 -4160 7190 -3970
rect -590 -4200 7190 -4160
rect 7810 -830 8390 -810
rect 7810 -3970 7830 -830
rect 8370 -3970 8390 -830
rect 7810 -4160 8390 -3970
rect 9010 -830 9590 -720
rect 9010 -3970 9030 -830
rect 9570 -3970 9590 -830
rect 9010 -4030 9590 -3970
rect 10210 -720 12650 -680
rect 10210 -830 10790 -720
rect 12610 -770 12650 -720
rect 13460 -710 13540 -670
rect 13460 -750 13480 -710
rect 13520 -750 13540 -710
rect 13760 -680 13800 -560
rect 15280 -590 15320 -70
rect 17060 -90 17080 -50
rect 17120 -90 17140 -50
rect 17410 -40 17990 30
rect 18610 3170 19190 3480
rect 19720 3370 23400 3390
rect 19720 3330 19740 3370
rect 19780 3350 23400 3370
rect 19780 3330 19800 3350
rect 19720 3310 19800 3330
rect 21240 3290 21320 3310
rect 21240 3250 21260 3290
rect 21300 3250 21320 3290
rect 21240 3230 21320 3250
rect 22460 3290 22540 3310
rect 22460 3250 22480 3290
rect 22520 3250 22540 3290
rect 22460 3230 22540 3250
rect 18610 30 18630 3170
rect 19170 30 19190 3170
rect 18610 10 19190 30
rect 19810 3170 20390 3190
rect 19810 30 19830 3170
rect 20370 30 20390 3170
rect 19810 -40 20390 30
rect 21010 3170 21590 3230
rect 21010 30 21030 3170
rect 21570 30 21590 3170
rect 21010 10 21590 30
rect 22210 3190 22790 3230
rect 22210 3170 23390 3190
rect 22210 30 22230 3170
rect 22770 30 22830 3170
rect 23370 30 23390 3170
rect 22210 10 23390 30
rect 17410 -80 20390 -40
rect 17060 -130 17140 -90
rect 17060 -170 17080 -130
rect 17120 -170 17140 -130
rect 17060 -190 17140 -170
rect 15280 -630 16790 -590
rect 13760 -720 15590 -680
rect 13460 -770 13540 -750
rect 10210 -3970 10230 -830
rect 10770 -3970 10790 -830
rect 9260 -4050 9340 -4030
rect 9260 -4090 9280 -4050
rect 9320 -4090 9340 -4050
rect 9260 -4110 9340 -4090
rect 10210 -4160 10790 -3970
rect 11410 -830 11990 -810
rect 11410 -3970 11430 -830
rect 11970 -3970 11990 -830
rect 11410 -4030 11990 -3970
rect 12610 -830 13190 -770
rect 12610 -3970 12630 -830
rect 13170 -3970 13190 -830
rect 12610 -3990 13190 -3970
rect 13810 -830 14390 -810
rect 13810 -3970 13830 -830
rect 14370 -3970 14390 -830
rect 7810 -4200 10790 -4160
rect 1070 -4690 1150 -4670
rect 1070 -4730 1090 -4690
rect 1130 -4710 1150 -4690
rect 1130 -4730 5990 -4710
rect 1070 -4750 5990 -4730
rect -3590 -4830 -2410 -4810
rect -3590 -7970 -3570 -4830
rect -3030 -7970 -2970 -4830
rect -2430 -7970 -2410 -4830
rect -3590 -7990 -2410 -7970
rect -2990 -8030 -2410 -7990
rect -1790 -4830 -1210 -4810
rect -1790 -7970 -1770 -4830
rect -1230 -7970 -1210 -4830
rect -1790 -8030 -1210 -7970
rect -590 -4830 -10 -4810
rect -590 -7970 -570 -4830
rect -30 -7970 -10 -4830
rect -590 -8030 -10 -7970
rect 610 -4830 1190 -4810
rect 610 -7970 630 -4830
rect 1170 -7970 1190 -4830
rect 610 -8030 1190 -7970
rect 1810 -4830 2990 -4810
rect 1810 -7970 1830 -4830
rect 2370 -7970 2430 -4830
rect 2970 -7970 2990 -4830
rect 1810 -7990 2990 -7970
rect 5410 -4830 5990 -4750
rect 6880 -4770 6920 -4200
rect 9260 -4710 9340 -4690
rect 9260 -4750 9280 -4710
rect 9320 -4750 9340 -4710
rect 9260 -4770 9340 -4750
rect 10480 -4770 10520 -4200
rect 11950 -4630 11990 -4030
rect 13810 -4160 14390 -3970
rect 15010 -830 15590 -720
rect 15010 -3970 15030 -830
rect 15570 -3970 15590 -830
rect 15010 -4030 15590 -3970
rect 16210 -830 16790 -630
rect 17680 -780 17720 -80
rect 20060 -710 20140 -690
rect 20060 -750 20080 -710
rect 20120 -750 20140 -710
rect 20060 -770 20140 -750
rect 21260 -710 21340 -690
rect 21260 -750 21280 -710
rect 21320 -750 21340 -710
rect 21260 -770 21340 -750
rect 22460 -710 22540 -690
rect 22460 -750 22480 -710
rect 22520 -750 22540 -710
rect 22460 -770 22540 -750
rect 16210 -3970 16230 -830
rect 16770 -3970 16790 -830
rect 15050 -4050 15130 -4030
rect 15050 -4090 15070 -4050
rect 15110 -4090 15130 -4050
rect 15050 -4110 15130 -4090
rect 16210 -4160 16790 -3970
rect 17410 -830 17990 -780
rect 17410 -3970 17430 -830
rect 17970 -3970 17990 -830
rect 17410 -4030 17990 -3970
rect 18610 -830 19190 -810
rect 18610 -3970 18630 -830
rect 19170 -3970 19190 -830
rect 17450 -4050 17530 -4030
rect 17450 -4090 17470 -4050
rect 17510 -4090 17530 -4050
rect 17450 -4110 17530 -4090
rect 18610 -4160 19190 -3970
rect 19810 -830 20390 -770
rect 19810 -3970 19830 -830
rect 20370 -3970 20390 -830
rect 19810 -3990 20390 -3970
rect 21010 -830 21590 -770
rect 21010 -3970 21030 -830
rect 21570 -3970 21590 -830
rect 21010 -3990 21590 -3970
rect 22210 -810 22790 -770
rect 22210 -830 23390 -810
rect 22210 -3970 22230 -830
rect 22770 -3970 22830 -830
rect 23370 -3970 23390 -830
rect 22210 -3990 23390 -3970
rect 13810 -4200 19190 -4160
rect 15050 -4610 15130 -4590
rect 15050 -4630 15070 -4610
rect 11950 -4650 15070 -4630
rect 15110 -4650 15130 -4610
rect 11950 -4670 15130 -4650
rect 5410 -7970 5430 -4830
rect 5970 -7970 5990 -4830
rect 5410 -7990 5990 -7970
rect 6610 -4830 7190 -4770
rect 6610 -7970 6630 -4830
rect 7170 -7970 7190 -4830
rect 6610 -7990 7190 -7970
rect 7810 -4830 8390 -4810
rect 7810 -7970 7830 -4830
rect 8370 -7970 8390 -4830
rect 7810 -7990 8390 -7970
rect 9010 -4830 9590 -4770
rect 9010 -7970 9030 -4830
rect 9570 -7970 9590 -4830
rect 9010 -7990 9590 -7970
rect 10210 -4830 10790 -4770
rect 10210 -7970 10230 -4830
rect 10770 -7970 10790 -4830
rect 10210 -7990 10790 -7970
rect 11410 -4830 11990 -4810
rect 11410 -7970 11430 -4830
rect 11970 -7970 11990 -4830
rect 11410 -7990 11990 -7970
rect 12610 -4830 13190 -4670
rect 15180 -4720 15220 -4200
rect 17450 -4700 17530 -4680
rect 17450 -4720 17470 -4700
rect 12610 -7970 12630 -4830
rect 13170 -7970 13190 -4830
rect 12610 -7990 13190 -7970
rect 13810 -4760 15220 -4720
rect 16210 -4740 17470 -4720
rect 17510 -4740 17530 -4700
rect 16210 -4760 17530 -4740
rect 13810 -4830 14390 -4760
rect 13810 -7970 13830 -4830
rect 14370 -7970 14390 -4830
rect 13810 -7990 14390 -7970
rect 15010 -4830 15590 -4810
rect 15010 -7970 15030 -4830
rect 15570 -7970 15590 -4830
rect 15010 -7990 15590 -7970
rect 16210 -4830 16790 -4760
rect 16210 -7970 16230 -4830
rect 16770 -7970 16790 -4830
rect 16210 -7990 16790 -7970
rect 17410 -4830 17990 -4810
rect 17410 -7970 17430 -4830
rect 17970 -7970 17990 -4830
rect 17410 -8030 17990 -7970
rect 18610 -4830 19190 -4810
rect 18610 -7970 18630 -4830
rect 19170 -7970 19190 -4830
rect 18610 -8030 19190 -7970
rect 19810 -4830 20390 -4810
rect 19810 -7970 19830 -4830
rect 20370 -7970 20390 -4830
rect 19810 -8030 20390 -7970
rect 21010 -4830 21590 -4810
rect 21010 -7970 21030 -4830
rect 21570 -7970 21590 -4830
rect 21010 -8030 21590 -7970
rect 22210 -4830 23390 -4810
rect 22210 -7970 22230 -4830
rect 22770 -7970 22830 -4830
rect 23370 -7970 23390 -4830
rect 22210 -7990 23390 -7970
rect 22210 -8030 22790 -7990
rect -2740 -8050 -2660 -8030
rect -2740 -8090 -2720 -8050
rect -2680 -8090 -2660 -8050
rect -2740 -8110 -2660 -8090
rect -1540 -8050 -1460 -8030
rect -1540 -8090 -1520 -8050
rect -1480 -8090 -1460 -8050
rect -1540 -8110 -1460 -8090
rect -340 -8050 -260 -8030
rect -340 -8090 -320 -8050
rect -280 -8090 -260 -8050
rect -340 -8110 -260 -8090
rect 860 -8050 940 -8030
rect 860 -8090 880 -8050
rect 920 -8090 940 -8050
rect 860 -8110 940 -8090
rect 6260 -8050 6340 -8030
rect 6260 -8090 6280 -8050
rect 6320 -8090 6340 -8050
rect 6260 -8180 6340 -8090
rect 6260 -8220 6280 -8180
rect 6320 -8220 6340 -8180
rect 7460 -8050 7540 -8030
rect 7460 -8090 7480 -8050
rect 7520 -8090 7540 -8050
rect 7460 -8130 7540 -8090
rect 7460 -8170 7480 -8130
rect 7520 -8170 7540 -8130
rect 7460 -8190 7540 -8170
rect 8660 -8050 8740 -8030
rect 8660 -8090 8680 -8050
rect 8720 -8090 8740 -8050
rect 8660 -8180 8740 -8090
rect 6260 -8240 6340 -8220
rect 8660 -8220 8680 -8180
rect 8720 -8220 8740 -8180
rect 8660 -8240 8740 -8220
rect 9860 -8050 9940 -8030
rect 9860 -8090 9880 -8050
rect 9920 -8090 9940 -8050
rect 9860 -8180 9940 -8090
rect 9860 -8220 9880 -8180
rect 9920 -8220 9940 -8180
rect 9860 -8240 9940 -8220
rect 11060 -8050 11140 -8030
rect 11060 -8090 11080 -8050
rect 11120 -8090 11140 -8050
rect 11060 -8180 11140 -8090
rect 11060 -8220 11080 -8180
rect 11120 -8220 11140 -8180
rect 11060 -8240 11140 -8220
rect 12260 -8050 12340 -8030
rect 12260 -8090 12280 -8050
rect 12320 -8090 12340 -8050
rect 12260 -8180 12340 -8090
rect 12260 -8220 12280 -8180
rect 12320 -8220 12340 -8180
rect 12260 -8240 12340 -8220
rect 13460 -8050 13540 -8030
rect 13460 -8090 13480 -8050
rect 13520 -8090 13540 -8050
rect 13460 -8180 13540 -8090
rect 13460 -8220 13480 -8180
rect 13520 -8220 13540 -8180
rect 13460 -8240 13540 -8220
rect 14660 -8050 14740 -8030
rect 14660 -8090 14680 -8050
rect 14720 -8090 14740 -8050
rect 14660 -8180 14740 -8090
rect 14660 -8220 14680 -8180
rect 14720 -8220 14740 -8180
rect 14660 -8240 14740 -8220
rect 15860 -8050 15940 -8030
rect 15860 -8090 15880 -8050
rect 15920 -8090 15940 -8050
rect 15860 -8180 15940 -8090
rect 17660 -8050 17740 -8030
rect 17660 -8090 17680 -8050
rect 17720 -8090 17740 -8050
rect 17660 -8110 17740 -8090
rect 18860 -8050 18940 -8030
rect 18860 -8090 18880 -8050
rect 18920 -8090 18940 -8050
rect 18860 -8110 18940 -8090
rect 20060 -8050 20140 -8030
rect 20060 -8090 20080 -8050
rect 20120 -8090 20140 -8050
rect 20060 -8110 20140 -8090
rect 21260 -8050 21340 -8030
rect 21260 -8090 21280 -8050
rect 21320 -8090 21340 -8050
rect 21260 -8110 21340 -8090
rect 22460 -8050 22540 -8030
rect 22460 -8090 22480 -8050
rect 22520 -8090 22540 -8050
rect 22460 -8110 22540 -8090
rect 15860 -8220 15880 -8180
rect 15920 -8220 15940 -8180
rect 15860 -8240 15940 -8220
<< viali >>
rect -3570 30 -3030 3170
rect -2970 30 -2430 3170
rect -1770 30 -1230 3170
rect 630 30 1170 3170
rect 6630 30 7170 3170
rect 7830 30 8370 3170
rect 5080 -170 5120 -130
rect 7480 -170 7520 -130
rect -3570 -3970 -3030 -830
rect -2970 -3970 -2430 -830
rect -1770 -3970 -1230 -830
rect 7480 -670 7520 -630
rect 11430 30 11970 3170
rect 9880 -170 9920 -130
rect 13830 30 14370 3170
rect 12280 -170 12320 -130
rect 16230 30 16770 3170
rect 14680 -170 14720 -130
rect 13480 -670 13520 -630
rect 21030 30 21570 3170
rect 22230 30 22770 3170
rect 22830 30 23370 3170
rect 17080 -170 17120 -130
rect -3570 -7970 -3030 -4830
rect -2970 -7970 -2430 -4830
rect -1770 -7970 -1230 -4830
rect -570 -7970 -30 -4830
rect 630 -7970 1170 -4830
rect 1830 -7970 2370 -4830
rect 19830 -3970 20370 -830
rect 21030 -3970 21570 -830
rect 22230 -3970 22770 -830
rect 22830 -3970 23370 -830
rect 7830 -7970 8370 -4830
rect 11430 -7970 11970 -4830
rect 15030 -7970 15570 -4830
rect 17430 -7970 17970 -4830
rect 18630 -7970 19170 -4830
rect 19830 -7970 20370 -4830
rect 21030 -7970 21570 -4830
rect 22230 -7970 22770 -4830
rect 22830 -7970 23370 -4830
rect 6280 -8220 6320 -8180
rect 7480 -8170 7520 -8130
rect 8680 -8220 8720 -8180
rect 9880 -8220 9920 -8180
rect 11080 -8220 11120 -8180
rect 12280 -8220 12320 -8180
rect 13480 -8220 13520 -8180
rect 14680 -8220 14720 -8180
rect 15880 -8220 15920 -8180
<< metal1 >>
rect -3600 3630 23400 6810
rect -3600 3170 -1210 3190
rect -3600 30 -3570 3170
rect -3030 30 -2970 3170
rect -2430 30 -1770 3170
rect -1230 30 -1210 3170
rect -3600 -800 -1210 30
rect 610 3170 1190 3630
rect 610 30 630 3170
rect 1170 30 1190 3170
rect 610 10 1190 30
rect 6610 3170 7190 3630
rect 6610 30 6630 3170
rect 7170 30 7190 3170
rect 6610 10 7190 30
rect 7810 3170 8390 3630
rect 7810 30 7830 3170
rect 8370 30 8390 3170
rect 7810 10 8390 30
rect 11410 3170 11990 3630
rect 11410 30 11430 3170
rect 11970 30 11990 3170
rect 11410 10 11990 30
rect 13810 3170 14390 3630
rect 13810 30 13830 3170
rect 14370 30 14390 3170
rect 13810 10 14390 30
rect 16210 3170 16790 3630
rect 16210 30 16230 3170
rect 16770 30 16790 3170
rect 16210 10 16790 30
rect 21010 3170 23390 3190
rect 21010 30 21030 3170
rect 21570 30 22230 3170
rect 22770 30 22830 3170
rect 23370 30 23390 3170
rect 5060 -130 5140 -110
rect 5060 -170 5080 -130
rect 5120 -170 5140 -130
rect 5060 -800 5140 -170
rect 7460 -130 7540 -30
rect 7460 -170 7480 -130
rect 7520 -170 7540 -130
rect 7460 -630 7540 -170
rect 7460 -670 7480 -630
rect 7520 -670 7540 -630
rect 7460 -800 7540 -670
rect 9860 -130 9940 -30
rect 9860 -170 9880 -130
rect 9920 -170 9940 -130
rect 9860 -800 9940 -170
rect 12260 -130 12340 -30
rect 12260 -170 12280 -130
rect 12320 -170 12340 -130
rect 12260 -800 12340 -170
rect 14660 -130 14740 -30
rect 14660 -170 14680 -130
rect 14720 -170 14740 -130
rect 13460 -630 13540 -610
rect 13460 -670 13480 -630
rect 13520 -670 13540 -630
rect 13460 -800 13540 -670
rect 14660 -800 14740 -170
rect 17060 -130 17140 -30
rect 17060 -170 17080 -130
rect 17120 -170 17140 -130
rect 17060 -800 17140 -170
rect 21010 -800 23390 30
rect -3600 -830 23400 -800
rect -3600 -3970 -3570 -830
rect -3030 -3970 -2970 -830
rect -2430 -3970 -1770 -830
rect -1230 -3970 19830 -830
rect 20370 -3970 21030 -830
rect 21570 -3970 22230 -830
rect 22770 -3970 22830 -830
rect 23370 -3970 23400 -830
rect -3600 -4830 23400 -3970
rect -3600 -7970 -3570 -4830
rect -3030 -7970 -2970 -4830
rect -2430 -7970 -1770 -4830
rect -1230 -7970 -570 -4830
rect -30 -7970 630 -4830
rect 1170 -7970 1830 -4830
rect 2370 -7970 7830 -4830
rect 8370 -7970 11430 -4830
rect 11970 -7970 15030 -4830
rect 15570 -7970 17430 -4830
rect 17970 -7970 18630 -4830
rect 19170 -7970 19830 -4830
rect 20370 -7970 21030 -4830
rect 21570 -7970 22230 -4830
rect 22770 -7970 22830 -4830
rect 23370 -7970 23400 -4830
rect -3600 -7990 23400 -7970
rect 6260 -8180 6340 -7990
rect 6260 -8220 6280 -8180
rect 6320 -8220 6340 -8180
rect 7460 -8130 7540 -7990
rect 7460 -8170 7480 -8130
rect 7520 -8170 7540 -8130
rect 7460 -8190 7540 -8170
rect 8660 -8180 8740 -7990
rect 6260 -8240 6340 -8220
rect 8660 -8220 8680 -8180
rect 8720 -8220 8740 -8180
rect 8660 -8240 8740 -8220
rect 9860 -8180 9940 -7990
rect 9860 -8220 9880 -8180
rect 9920 -8220 9940 -8180
rect 9860 -8240 9940 -8220
rect 11060 -8180 11140 -7990
rect 11060 -8220 11080 -8180
rect 11120 -8220 11140 -8180
rect 11060 -8240 11140 -8220
rect 12260 -8180 12340 -7990
rect 12260 -8220 12280 -8180
rect 12320 -8220 12340 -8180
rect 12260 -8240 12340 -8220
rect 13460 -8180 13540 -7990
rect 13460 -8220 13480 -8180
rect 13520 -8220 13540 -8180
rect 13460 -8240 13540 -8220
rect 14660 -8180 14740 -7990
rect 14660 -8220 14680 -8180
rect 14720 -8220 14740 -8180
rect 14660 -8240 14740 -8220
rect 15860 -8180 15940 -7990
rect 15860 -8220 15880 -8180
rect 15920 -8220 15940 -8180
rect 15860 -8240 15940 -8220
<< end >>
