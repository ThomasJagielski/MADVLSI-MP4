magic
tech sky130A
timestamp 1617673688
<< nwell >>
rect 7125 1060 7515 1120
<< nmos >>
rect 3530 -6525 3930 -6520
rect 4330 -6525 4730 -6520
rect 5930 -6525 6330 -6520
rect 6730 -6525 7130 -6520
rect 8330 -6525 8730 -6520
rect 9130 -6525 9530 -6520
<< ndiffc >>
rect -14925 -5245 -14905 -5175
rect -13325 -5245 -13305 -5175
rect -12525 -5245 -12505 -5175
rect -10925 -5245 -10905 -5175
rect -10125 -5245 -10105 -5175
rect -8525 -5245 -8505 -5175
rect -7725 -5245 -7705 -5175
<< poly >>
rect 7125 1105 7515 1115
rect 7125 1085 7135 1105
rect 7505 1085 7515 1105
rect 7125 925 7515 1085
rect 7125 905 7135 925
rect 7505 905 7515 925
rect 7125 895 7515 905
rect 3530 -6560 3930 -6525
rect 3530 -6580 3540 -6560
rect 3920 -6580 3930 -6560
rect 3530 -6590 3930 -6580
rect 4330 -6560 4730 -6525
rect 4330 -6580 4340 -6560
rect 4720 -6580 4730 -6560
rect 4330 -6590 4730 -6580
rect 5930 -6560 6330 -6525
rect 5930 -6580 5940 -6560
rect 6320 -6580 6330 -6560
rect 5930 -6590 6330 -6580
rect 6730 -6560 7130 -6525
rect 6730 -6580 6740 -6560
rect 7120 -6580 7130 -6560
rect 6730 -6590 7130 -6580
rect 8330 -6560 8730 -6525
rect 8330 -6580 8340 -6560
rect 8720 -6580 8730 -6560
rect 8330 -6590 8730 -6580
rect 9130 -6560 9530 -6525
rect 9130 -6580 9140 -6560
rect 9520 -6580 9530 -6560
rect 9130 -6590 9530 -6580
<< polycont >>
rect 7135 1085 7505 1105
rect 7135 905 7505 925
rect 3540 -6580 3920 -6560
rect 4340 -6580 4720 -6560
rect 5940 -6580 6320 -6560
rect 6740 -6580 7120 -6560
rect 8340 -6580 8720 -6560
rect 9140 -6580 9520 -6560
<< locali >>
rect -2775 1230 -2125 1270
rect -2165 1040 -2125 1230
rect 7125 1105 7515 1180
rect 7125 1085 7135 1105
rect 7505 1085 7515 1105
rect 7125 1075 7515 1085
rect -2165 1020 -2100 1040
rect 9545 1000 9915 1175
rect 9545 960 11525 1000
rect 7125 925 9925 935
rect 7125 905 7135 925
rect 7505 905 9925 925
rect 7125 895 9925 905
rect 9535 -930 9925 895
rect 11135 -745 11525 960
rect -19825 -2760 -19370 -2660
rect -19470 -5490 -19370 -2760
rect -13380 -4540 -13360 -4535
rect -15000 -4835 -14960 -4575
rect -13400 -4835 -13360 -4540
rect -12600 -4835 -12560 -4535
rect -11000 -4835 -10960 -4560
rect -10200 -4835 -10160 -4570
rect -8600 -4835 -8560 -4570
rect -7800 -4835 -7760 -4570
rect -15370 -5295 -15185 -5275
rect -13770 -5295 -13685 -5275
rect -12970 -5295 -12885 -5275
rect -11370 -5295 -11285 -5275
rect -10570 -5295 -10485 -5275
rect -8970 -5295 -8885 -5275
rect -8170 -5295 -8085 -5275
rect -15370 -5490 -15345 -5295
rect -13770 -5490 -13745 -5295
rect -12970 -5490 -12945 -5295
rect -11370 -5490 -11345 -5295
rect -10570 -5490 -10545 -5295
rect -8970 -5490 -8945 -5295
rect -8170 -5490 -8145 -5295
rect -19470 -5590 -2710 -5490
rect -2810 -6740 -2710 -5590
rect 1930 -6740 2330 -6550
rect 3530 -6560 3930 -6550
rect 3530 -6580 3540 -6560
rect 3920 -6580 3930 -6560
rect 3530 -6590 3930 -6580
rect 4330 -6560 4730 -6550
rect 4330 -6580 4340 -6560
rect 4720 -6580 4730 -6560
rect 4330 -6590 4730 -6580
rect 5930 -6560 6330 -6550
rect 5930 -6580 5940 -6560
rect 6320 -6580 6330 -6560
rect 5930 -6590 6330 -6580
rect 6730 -6560 7130 -6550
rect 6730 -6580 6740 -6560
rect 7120 -6580 7130 -6560
rect 6730 -6590 7130 -6580
rect 8330 -6560 8730 -6550
rect 8330 -6580 8340 -6560
rect 8720 -6580 8730 -6560
rect 8330 -6590 8730 -6580
rect 9130 -6560 9530 -6550
rect 9130 -6580 9140 -6560
rect 9520 -6580 9530 -6560
rect 9130 -6590 9530 -6580
rect -2810 -6840 2330 -6740
<< viali >>
rect -14925 -5245 -14905 -5175
rect -13325 -5245 -13305 -5175
rect -12525 -5245 -12505 -5175
rect -10925 -5245 -10905 -5175
rect -10125 -5245 -10105 -5175
rect -8525 -5245 -8505 -5175
rect -7725 -5245 -7705 -5175
rect 3540 -6580 3920 -6560
rect 4340 -6580 4720 -6560
rect 5940 -6580 6320 -6560
rect 6740 -6580 7120 -6560
rect 8340 -6580 8720 -6560
rect 9140 -6580 9520 -6560
<< metal1 >>
rect -19820 1940 -18975 2895
rect -11975 1380 -11575 1385
rect -11975 1310 -11970 1380
rect -11580 1310 -11575 1380
rect -11975 1305 -11575 1310
rect -2935 1300 14320 2895
rect -2070 -295 14320 1300
rect -15285 -4945 -7670 -4830
rect -15285 -5015 -11970 -4945
rect -11580 -5015 -7670 -4945
rect -15285 -5020 -7670 -5015
rect -15285 -5175 -14870 -5100
rect -15285 -5245 -14925 -5175
rect -14905 -5245 -14870 -5175
rect -15285 -5455 -14870 -5245
rect -13685 -5175 -13270 -5075
rect -13685 -5245 -13325 -5175
rect -13305 -5245 -13270 -5175
rect -13685 -5455 -13270 -5245
rect -12885 -5175 -12470 -5115
rect -12885 -5245 -12525 -5175
rect -12505 -5245 -12470 -5175
rect -12885 -5455 -12470 -5245
rect -11285 -5175 -10870 -5085
rect -11285 -5245 -10925 -5175
rect -10905 -5245 -10870 -5175
rect -11285 -5455 -10870 -5245
rect -10485 -5175 -10070 -5090
rect -10485 -5245 -10125 -5175
rect -10105 -5245 -10070 -5175
rect -10485 -5455 -10070 -5245
rect -8885 -5175 -8470 -5085
rect -8885 -5245 -8525 -5175
rect -8505 -5245 -8470 -5175
rect -8885 -5455 -8470 -5245
rect -8085 -5175 -7670 -5105
rect -8085 -5245 -7725 -5175
rect -7705 -5245 -7670 -5175
rect -8085 -5455 -7670 -5245
rect -20905 -6560 14330 -5455
rect -20905 -6580 3540 -6560
rect 3920 -6580 4340 -6560
rect 4720 -6580 5940 -6560
rect 6320 -6580 6740 -6560
rect 7120 -6580 8340 -6560
rect 8720 -6580 9140 -6560
rect 9520 -6580 14330 -6560
rect -20905 -8000 14330 -6580
<< via1 >>
rect -11970 1310 -11580 1380
rect -11970 -5015 -11580 -4945
<< metal2 >>
rect -11975 1380 -11575 1385
rect -11975 1310 -11970 1380
rect -11580 1310 -11575 1380
rect -11975 -4945 -11575 1310
rect -11975 -5015 -11970 -4945
rect -11580 -5015 -11575 -4945
rect -11975 -5020 -11575 -5015
use low-voltage_super-wilson  low-voltage_super-wilson_0
timestamp 1617673688
transform 1 0 -1485 0 1 1175
box -615 -275 15825 1785
use mux2  mux2_0
timestamp 1617673688
transform 1 0 -15285 0 1 -5275
box 0 -60 415 505
use mux2  mux2_1
timestamp 1617673688
transform 1 0 -13685 0 1 -5275
box 0 -60 415 505
use mux2  mux2_2
timestamp 1617673688
transform 1 0 -12885 0 1 -5275
box 0 -60 415 505
use mux2  mux2_3
timestamp 1617673688
transform 1 0 -11285 0 1 -5275
box 0 -60 415 505
use mux2  mux2_4
timestamp 1617673688
transform 1 0 -10485 0 1 -5275
box 0 -60 415 505
use mux2  mux2_5
timestamp 1617673688
transform 1 0 -8885 0 1 -5275
box 0 -60 415 505
use mux2  mux2_6
timestamp 1617673688
transform 1 0 -8085 0 1 -5275
box 0 -60 415 505
use dac_ladder  dac_ladder_0
timestamp 1617673688
transform 1 0 2630 0 1 -2525
box -4700 -4135 11700 3405
use dac_ladder  dac_ladder_1
timestamp 1617673688
transform 1 0 -14475 0 1 -510
box -4700 -4135 11700 3405
use ibias_vg  ibias_vg_0
timestamp 1617673688
transform 1 0 -43680 0 1 300
box -820 -8300 24030 2600
<< labels >>
rlabel poly 3785 -6590 3785 -6590 5 b0
rlabel poly 4585 -6590 4585 -6590 5 b0
rlabel poly 6185 -6590 6185 -6590 5 b0
rlabel poly 6985 -6590 6985 -6590 5 b0
rlabel poly 8585 -6590 8585 -6590 5 b0
rlabel poly 9385 -6590 9385 -6590 5 b0
rlabel metal1 -13685 -5325 -13685 -5325 7 B
rlabel locali -13685 -5285 -13685 -5285 7 A
rlabel locali -12885 -5285 -12885 -5285 7 A
rlabel metal1 -12885 -5325 -12885 -5325 7 B
rlabel metal1 -11285 -5325 -11285 -5325 7 B
rlabel locali -11285 -5285 -11285 -5285 7 A
rlabel metal1 -10485 -5325 -10485 -5325 7 B
rlabel locali -10485 -5285 -10485 -5285 7 A
rlabel metal1 -8885 -5325 -8885 -5325 7 B
rlabel locali -8885 -5285 -8885 -5285 7 A
rlabel locali -8085 -5285 -8085 -5285 7 A
rlabel metal1 -8085 -5325 -8085 -5325 7 B
<< end >>
