magic
tech sky130A
magscale 1 2
timestamp 1617377580
<< error_p >>
rect 2400 10 3200 3210
rect 10738 2060 10830 2512
rect 10738 10 11200 2060
rect 12000 10 12800 2060
rect 13600 10 14400 1980
rect 15200 10 16000 1980
rect 16800 10 17600 2512
rect 18400 10 19200 2512
rect 2400 -4790 3200 -1590
rect 4000 -4790 4800 -2428
rect 5600 -4790 6400 -2820
rect 7200 -4790 8000 -2820
rect 8800 -4790 9600 -2820
rect 10400 -4790 11200 -2820
rect 12000 -4790 12800 -2820
rect 13600 -4790 14400 -2820
rect 15200 -4790 16000 -2820
rect 16800 -4790 17600 -1590
rect 18400 -4790 19200 -1590
rect 20000 -3687 20800 -2933
rect 2400 -9830 3200 -6630
rect 4000 -9830 4800 -6630
rect 5600 -9830 6400 -6630
rect 7200 -9830 8000 -7860
rect 8800 -9830 9600 -7860
rect 10400 -9830 11200 -7860
rect 12000 -9830 12800 -7860
rect 13600 -9830 14400 -7860
rect 15200 -9830 16000 -7860
rect 16800 -9830 17600 -7860
rect 18400 -9830 19200 -6630
rect 2400 -14630 3200 -11430
rect 4000 -14630 4800 -11430
rect 5600 -13130 6400 -11430
rect 7200 -13130 8000 -11430
rect 8800 -13130 9600 -11430
rect 10400 -14630 11200 -11430
rect 12000 -14630 12800 -11430
rect 13600 -13400 14400 -11430
rect 15200 -13400 16000 -11430
rect 16800 -13400 17600 -11430
rect 18400 -13400 18740 -11430
<< nmos >>
rect 0 10 800 3210
rect 1600 10 2400 3210
rect 3200 10 4000 3210
rect 4800 10 5600 3210
rect 6400 10 7200 3210
rect 8000 10 8800 3210
rect 9600 10 10400 3210
rect 11200 10 12000 3210
rect 12800 10 13600 3210
rect 14400 10 15200 3210
rect 16000 10 16800 3210
rect 17600 10 18400 3210
rect 19200 10 20000 3210
rect 20800 10 21600 3210
rect 24000 10 24800 3210
rect 25600 10 26400 3210
rect 27200 10 28000 3210
rect 28800 10 29600 3210
rect 30400 10 31200 3210
rect 32000 10 32800 3210
rect 37600 10 38400 3210
rect 39200 10 40000 3210
rect 40800 10 41600 3210
rect 42400 10 43200 3210
rect 44000 10 44800 3210
rect 45600 10 46400 3210
rect 0 -4790 800 -1590
rect 1600 -4790 2400 -1590
rect 3200 -4790 4000 -1590
rect 4800 -4790 5600 -1590
rect 6400 -4790 7200 -1590
rect 8000 -4790 8800 -1590
rect 9600 -4790 10400 -1590
rect 11200 -4790 12000 -1590
rect 12800 -4790 13600 -1590
rect 14400 -4790 15200 -1590
rect 16000 -4790 16800 -1590
rect 17600 -4790 18400 -1590
rect 19200 -4790 20000 -1590
rect 20800 -4790 21600 -1590
rect 24000 -4790 24800 -1590
rect 25600 -4790 26400 -1590
rect 27200 -4790 28000 -1590
rect 28800 -4790 29600 -1590
rect 30400 -4790 31200 -1590
rect 32000 -4790 32800 -1590
rect 37600 -4790 38400 -1590
rect 39200 -4790 40000 -1590
rect 40800 -4790 41600 -1590
rect 42400 -4790 43200 -1590
rect 44000 -4790 44800 -1590
rect 45600 -4790 46400 -1590
rect 0 -9830 800 -6630
rect 1600 -9830 2400 -6630
rect 3200 -9830 4000 -6630
rect 4800 -9830 5600 -6630
rect 6400 -9830 7200 -6630
rect 8000 -9830 8800 -6630
rect 9600 -9830 10400 -6630
rect 11200 -9830 12000 -6630
rect 12800 -9830 13600 -6630
rect 14400 -9830 15200 -6630
rect 16000 -9830 16800 -6630
rect 17600 -9830 18400 -6630
rect 19200 -9830 20000 -6630
rect 20800 -9830 21600 -6630
rect 24000 -9830 24800 -6630
rect 25600 -9830 26400 -6630
rect 27200 -9830 28000 -6630
rect 28800 -9830 29600 -6630
rect 30400 -9830 31200 -6630
rect 32000 -9830 32800 -6630
rect 37600 -9830 38400 -6630
rect 39200 -9830 40000 -6630
rect 40800 -9830 41600 -6630
rect 42400 -9830 43200 -6630
rect 44000 -9830 44800 -6630
rect 45600 -9830 46400 -6630
rect 0 -14630 800 -11430
rect 1600 -14630 2400 -11430
rect 3200 -14630 4000 -11430
rect 4800 -14630 5600 -11430
rect 6400 -14630 7200 -11430
rect 8000 -14630 8800 -11430
rect 9600 -14630 10400 -11430
rect 11200 -14630 12000 -11430
rect 12800 -14630 13600 -11430
rect 14400 -14630 15200 -11430
rect 16000 -14630 16800 -11430
rect 17600 -14630 18400 -11430
rect 19200 -14630 20000 -11430
rect 20800 -14630 21600 -11430
rect 24000 -14630 24800 -11430
rect 25600 -14630 26400 -11430
rect 27200 -14630 28000 -11430
rect 28800 -14630 29600 -11430
rect 30400 -14630 31200 -11430
rect 32000 -14630 32800 -11430
rect 37600 -14630 38400 -11430
rect 39200 -14630 40000 -11430
rect 40800 -14630 41600 -11430
rect 42400 -14630 43200 -11430
rect 44000 -14630 44800 -11430
rect 45600 -14630 46400 -11430
<< ndiff >>
rect -800 3170 0 3210
rect -800 50 -760 3170
rect -40 50 0 3170
rect -800 10 0 50
rect 800 3170 1600 3210
rect 800 50 840 3170
rect 1560 50 1600 3170
rect 800 10 1600 50
rect 2400 3170 3200 3210
rect 2400 50 2440 3170
rect 3160 50 3200 3170
rect 2400 10 3200 50
rect 4000 3170 4800 3210
rect 4000 50 4040 3170
rect 4760 50 4800 3170
rect 4000 10 4800 50
rect 5600 3170 6400 3210
rect 5600 50 5640 3170
rect 6360 50 6400 3170
rect 5600 10 6400 50
rect 7200 3170 8000 3210
rect 7200 50 7240 3170
rect 7960 50 8000 3170
rect 7200 10 8000 50
rect 8800 3170 9600 3210
rect 8800 50 8840 3170
rect 9560 50 9600 3170
rect 8800 10 9600 50
rect 10400 3170 11200 3210
rect 10400 50 10440 3170
rect 11160 50 11200 3170
rect 10400 10 11200 50
rect 12000 3170 12800 3210
rect 12000 50 12040 3170
rect 12760 50 12800 3170
rect 12000 10 12800 50
rect 13600 3170 14400 3210
rect 13600 50 13640 3170
rect 14360 50 14400 3170
rect 13600 10 14400 50
rect 15200 3170 16000 3210
rect 15200 50 15240 3170
rect 15960 50 16000 3170
rect 15200 10 16000 50
rect 16800 3170 17600 3210
rect 16800 50 16840 3170
rect 17560 50 17600 3170
rect 16800 10 17600 50
rect 18400 3170 19200 3210
rect 18400 50 18440 3170
rect 19160 50 19200 3170
rect 18400 10 19200 50
rect 20000 3170 20800 3210
rect 20000 50 20040 3170
rect 20760 50 20800 3170
rect 20000 10 20800 50
rect 21600 3170 22400 3210
rect 23200 3170 24000 3210
rect 21600 50 21640 3170
rect 22360 50 22400 3170
rect 23200 50 23240 3170
rect 23960 50 24000 3170
rect 21600 10 22400 50
rect 23200 10 24000 50
rect 24800 3170 25600 3210
rect 24800 50 24840 3170
rect 25560 50 25600 3170
rect 24800 10 25600 50
rect 26400 3170 27200 3210
rect 26400 50 26440 3170
rect 27160 50 27200 3170
rect 26400 10 27200 50
rect 28000 3170 28800 3210
rect 28000 50 28040 3170
rect 28760 50 28800 3170
rect 28000 10 28800 50
rect 29600 3170 30400 3210
rect 29600 50 29640 3170
rect 30360 50 30400 3170
rect 29600 10 30400 50
rect 31200 3170 32000 3210
rect 31200 50 31240 3170
rect 31960 50 32000 3170
rect 31200 10 32000 50
rect 32800 3170 33600 3210
rect 32800 50 32840 3170
rect 33560 50 33600 3170
rect 32800 10 33600 50
rect 36800 3170 37600 3210
rect 36800 50 36840 3170
rect 37560 50 37600 3170
rect 36800 10 37600 50
rect 38400 3170 39200 3210
rect 38400 50 38440 3170
rect 39160 50 39200 3170
rect 38400 10 39200 50
rect 40000 3170 40800 3210
rect 40000 50 40040 3170
rect 40760 50 40800 3170
rect 40000 10 40800 50
rect 41600 3170 42400 3210
rect 41600 50 41640 3170
rect 42360 50 42400 3170
rect 41600 10 42400 50
rect 43200 3170 44000 3210
rect 43200 50 43240 3170
rect 43960 50 44000 3170
rect 43200 10 44000 50
rect 44800 3170 45600 3210
rect 44800 50 44840 3170
rect 45560 50 45600 3170
rect 44800 10 45600 50
rect 46400 3170 47200 3210
rect 46400 50 46440 3170
rect 47160 50 47200 3170
rect 46400 10 47200 50
rect -800 -1630 0 -1590
rect -800 -4750 -760 -1630
rect -40 -4750 0 -1630
rect -800 -4790 0 -4750
rect 800 -1630 1600 -1590
rect 800 -4750 840 -1630
rect 1560 -4750 1600 -1630
rect 800 -4790 1600 -4750
rect 2400 -1630 3200 -1590
rect 2400 -4750 2440 -1630
rect 3160 -4750 3200 -1630
rect 2400 -4790 3200 -4750
rect 4000 -1630 4800 -1590
rect 4000 -4750 4040 -1630
rect 4760 -4750 4800 -1630
rect 4000 -4790 4800 -4750
rect 5600 -1630 6400 -1590
rect 5600 -4750 5640 -1630
rect 6360 -4750 6400 -1630
rect 5600 -4790 6400 -4750
rect 7200 -1630 8000 -1590
rect 7200 -4750 7240 -1630
rect 7960 -4750 8000 -1630
rect 7200 -4790 8000 -4750
rect 8800 -1630 9600 -1590
rect 8800 -4750 8840 -1630
rect 9560 -4750 9600 -1630
rect 8800 -4790 9600 -4750
rect 10400 -1630 11200 -1590
rect 10400 -4750 10440 -1630
rect 11160 -4750 11200 -1630
rect 10400 -4790 11200 -4750
rect 12000 -1630 12800 -1590
rect 12000 -4750 12040 -1630
rect 12760 -4750 12800 -1630
rect 12000 -4790 12800 -4750
rect 13600 -1630 14400 -1590
rect 13600 -4750 13640 -1630
rect 14360 -4750 14400 -1630
rect 13600 -4790 14400 -4750
rect 15200 -1630 16000 -1590
rect 15200 -4750 15240 -1630
rect 15960 -4750 16000 -1630
rect 15200 -4790 16000 -4750
rect 16800 -1630 17600 -1590
rect 16800 -4750 16840 -1630
rect 17560 -4750 17600 -1630
rect 16800 -4790 17600 -4750
rect 18400 -1630 19200 -1590
rect 18400 -4750 18440 -1630
rect 19160 -4750 19200 -1630
rect 18400 -4790 19200 -4750
rect 20000 -1630 20800 -1590
rect 20000 -4750 20040 -1630
rect 20760 -4750 20800 -1630
rect 20000 -4790 20800 -4750
rect 21600 -1630 22400 -1590
rect 23200 -1630 24000 -1590
rect 21600 -4750 21640 -1630
rect 22360 -4750 22400 -1630
rect 23200 -4750 23240 -1630
rect 23960 -4750 24000 -1630
rect 21600 -4790 22400 -4750
rect 23200 -4790 24000 -4750
rect 24800 -1630 25600 -1590
rect 24800 -4750 24840 -1630
rect 25560 -4750 25600 -1630
rect 24800 -4790 25600 -4750
rect 26400 -1630 27200 -1590
rect 26400 -4750 26440 -1630
rect 27160 -4750 27200 -1630
rect 26400 -4790 27200 -4750
rect 28000 -1630 28800 -1590
rect 28000 -4750 28040 -1630
rect 28760 -4750 28800 -1630
rect 28000 -4790 28800 -4750
rect 29600 -1630 30400 -1590
rect 29600 -4750 29640 -1630
rect 30360 -4750 30400 -1630
rect 29600 -4790 30400 -4750
rect 31200 -1630 32000 -1590
rect 31200 -4750 31240 -1630
rect 31960 -4750 32000 -1630
rect 31200 -4790 32000 -4750
rect 32800 -1630 33600 -1590
rect 32800 -4750 32840 -1630
rect 33560 -4750 33600 -1630
rect 32800 -4790 33600 -4750
rect 36800 -1630 37600 -1590
rect 36800 -4750 36840 -1630
rect 37560 -4750 37600 -1630
rect 36800 -4790 37600 -4750
rect 38400 -1630 39200 -1590
rect 38400 -4750 38440 -1630
rect 39160 -4750 39200 -1630
rect 38400 -4790 39200 -4750
rect 40000 -1630 40800 -1590
rect 40000 -4750 40040 -1630
rect 40760 -4750 40800 -1630
rect 40000 -4790 40800 -4750
rect 41600 -1630 42400 -1590
rect 41600 -4750 41640 -1630
rect 42360 -4750 42400 -1630
rect 41600 -4790 42400 -4750
rect 43200 -1630 44000 -1590
rect 43200 -4750 43240 -1630
rect 43960 -4750 44000 -1630
rect 43200 -4790 44000 -4750
rect 44800 -1630 45600 -1590
rect 44800 -4750 44840 -1630
rect 45560 -4750 45600 -1630
rect 44800 -4790 45600 -4750
rect 46400 -1630 47200 -1590
rect 46400 -4750 46440 -1630
rect 47160 -4750 47200 -1630
rect 46400 -4790 47200 -4750
rect -800 -6670 0 -6630
rect -800 -9790 -760 -6670
rect -40 -9790 0 -6670
rect -800 -9830 0 -9790
rect 800 -6670 1600 -6630
rect 800 -9790 840 -6670
rect 1560 -9790 1600 -6670
rect 800 -9830 1600 -9790
rect 2400 -6670 3200 -6630
rect 2400 -9790 2440 -6670
rect 3160 -9790 3200 -6670
rect 2400 -9830 3200 -9790
rect 4000 -6670 4800 -6630
rect 4000 -9790 4040 -6670
rect 4760 -9790 4800 -6670
rect 4000 -9830 4800 -9790
rect 5600 -6670 6400 -6630
rect 5600 -9790 5640 -6670
rect 6360 -9790 6400 -6670
rect 5600 -9830 6400 -9790
rect 7200 -6670 8000 -6630
rect 7200 -9790 7240 -6670
rect 7960 -9790 8000 -6670
rect 7200 -9830 8000 -9790
rect 8800 -6670 9600 -6630
rect 8800 -9790 8840 -6670
rect 9560 -9790 9600 -6670
rect 8800 -9830 9600 -9790
rect 10400 -6670 11200 -6630
rect 10400 -9790 10440 -6670
rect 11160 -9790 11200 -6670
rect 10400 -9830 11200 -9790
rect 12000 -6670 12800 -6630
rect 12000 -9790 12040 -6670
rect 12760 -9790 12800 -6670
rect 12000 -9830 12800 -9790
rect 13600 -6670 14400 -6630
rect 13600 -9790 13640 -6670
rect 14360 -9790 14400 -6670
rect 13600 -9830 14400 -9790
rect 15200 -6670 16000 -6630
rect 15200 -9790 15240 -6670
rect 15960 -9790 16000 -6670
rect 15200 -9830 16000 -9790
rect 16800 -6670 17600 -6630
rect 16800 -9790 16840 -6670
rect 17560 -9790 17600 -6670
rect 16800 -9830 17600 -9790
rect 18400 -6670 19200 -6630
rect 18400 -9790 18440 -6670
rect 19160 -9790 19200 -6670
rect 18400 -9830 19200 -9790
rect 20000 -6670 20800 -6630
rect 20000 -9790 20040 -6670
rect 20760 -9790 20800 -6670
rect 20000 -9830 20800 -9790
rect 21600 -6670 22400 -6630
rect 23200 -6670 24000 -6630
rect 21600 -9790 21640 -6670
rect 22360 -9790 22400 -6670
rect 23200 -9790 23240 -6670
rect 23960 -9790 24000 -6670
rect 21600 -9830 22400 -9790
rect 23200 -9830 24000 -9790
rect 24800 -6670 25600 -6630
rect 24800 -9790 24840 -6670
rect 25560 -9790 25600 -6670
rect 24800 -9830 25600 -9790
rect 26400 -6670 27200 -6630
rect 26400 -9790 26440 -6670
rect 27160 -9790 27200 -6670
rect 26400 -9830 27200 -9790
rect 28000 -6670 28800 -6630
rect 28000 -9790 28040 -6670
rect 28760 -9790 28800 -6670
rect 28000 -9830 28800 -9790
rect 29600 -6670 30400 -6630
rect 29600 -9790 29640 -6670
rect 30360 -9790 30400 -6670
rect 29600 -9830 30400 -9790
rect 31200 -6670 32000 -6630
rect 31200 -9790 31240 -6670
rect 31960 -9790 32000 -6670
rect 31200 -9830 32000 -9790
rect 32800 -6670 33600 -6630
rect 32800 -9790 32840 -6670
rect 33560 -9790 33600 -6670
rect 32800 -9830 33600 -9790
rect 36800 -6670 37600 -6630
rect 36800 -9790 36840 -6670
rect 37560 -9790 37600 -6670
rect 36800 -9830 37600 -9790
rect 38400 -6670 39200 -6630
rect 38400 -9790 38440 -6670
rect 39160 -9790 39200 -6670
rect 38400 -9830 39200 -9790
rect 40000 -6670 40800 -6630
rect 40000 -9790 40040 -6670
rect 40760 -9790 40800 -6670
rect 40000 -9830 40800 -9790
rect 41600 -6670 42400 -6630
rect 41600 -9790 41640 -6670
rect 42360 -9790 42400 -6670
rect 41600 -9830 42400 -9790
rect 43200 -6670 44000 -6630
rect 43200 -9790 43240 -6670
rect 43960 -9790 44000 -6670
rect 43200 -9830 44000 -9790
rect 44800 -6670 45600 -6630
rect 44800 -9790 44840 -6670
rect 45560 -9790 45600 -6670
rect 44800 -9830 45600 -9790
rect 46400 -6670 47200 -6630
rect 46400 -9790 46440 -6670
rect 47160 -9790 47200 -6670
rect 46400 -9830 47200 -9790
rect -800 -11470 0 -11430
rect -800 -14590 -760 -11470
rect -40 -14590 0 -11470
rect -800 -14630 0 -14590
rect 800 -11470 1600 -11430
rect 800 -14590 840 -11470
rect 1560 -14590 1600 -11470
rect 800 -14630 1600 -14590
rect 2400 -11470 3200 -11430
rect 2400 -14590 2440 -11470
rect 3160 -14590 3200 -11470
rect 2400 -14630 3200 -14590
rect 4000 -11470 4800 -11430
rect 4000 -14590 4040 -11470
rect 4760 -14590 4800 -11470
rect 4000 -14630 4800 -14590
rect 5600 -11470 6400 -11430
rect 5600 -14590 5640 -11470
rect 6360 -14590 6400 -11470
rect 5600 -14630 6400 -14590
rect 7200 -11470 8000 -11430
rect 7200 -14590 7240 -11470
rect 7960 -14590 8000 -11470
rect 7200 -14630 8000 -14590
rect 8800 -11470 9600 -11430
rect 8800 -14590 8840 -11470
rect 9560 -14590 9600 -11470
rect 8800 -14630 9600 -14590
rect 10400 -11470 11200 -11430
rect 10400 -14590 10440 -11470
rect 11160 -14590 11200 -11470
rect 10400 -14630 11200 -14590
rect 12000 -11470 12800 -11430
rect 12000 -14590 12040 -11470
rect 12760 -14590 12800 -11470
rect 12000 -14630 12800 -14590
rect 13600 -11470 14400 -11430
rect 13600 -14590 13640 -11470
rect 14360 -14590 14400 -11470
rect 13600 -14630 14400 -14590
rect 15200 -11470 16000 -11430
rect 15200 -14590 15240 -11470
rect 15960 -14590 16000 -11470
rect 15200 -14630 16000 -14590
rect 16800 -11470 17600 -11430
rect 16800 -14590 16840 -11470
rect 17560 -14590 17600 -11470
rect 16800 -14630 17600 -14590
rect 18400 -11470 19200 -11430
rect 18400 -14590 18440 -11470
rect 19160 -14590 19200 -11470
rect 18400 -14630 19200 -14590
rect 20000 -11470 20800 -11430
rect 20000 -14590 20040 -11470
rect 20760 -14590 20800 -11470
rect 20000 -14630 20800 -14590
rect 21600 -11470 22400 -11430
rect 23200 -11470 24000 -11430
rect 21600 -14590 21640 -11470
rect 22360 -14590 22400 -11470
rect 23200 -14590 23240 -11470
rect 23960 -14590 24000 -11470
rect 21600 -14630 22400 -14590
rect 23200 -14630 24000 -14590
rect 24800 -11470 25600 -11430
rect 24800 -14590 24840 -11470
rect 25560 -14590 25600 -11470
rect 24800 -14630 25600 -14590
rect 26400 -11470 27200 -11430
rect 26400 -14590 26440 -11470
rect 27160 -14590 27200 -11470
rect 26400 -14630 27200 -14590
rect 28000 -11470 28800 -11430
rect 28000 -14590 28040 -11470
rect 28760 -14590 28800 -11470
rect 28000 -14630 28800 -14590
rect 29600 -11470 30400 -11430
rect 29600 -14590 29640 -11470
rect 30360 -14590 30400 -11470
rect 29600 -14630 30400 -14590
rect 31200 -11470 32000 -11430
rect 31200 -14590 31240 -11470
rect 31960 -14590 32000 -11470
rect 31200 -14630 32000 -14590
rect 32800 -11470 33600 -11430
rect 32800 -14590 32840 -11470
rect 33560 -14590 33600 -11470
rect 32800 -14630 33600 -14590
rect 36800 -11470 37600 -11430
rect 36800 -14590 36840 -11470
rect 37560 -14590 37600 -11470
rect 36800 -14630 37600 -14590
rect 38400 -11470 39200 -11430
rect 38400 -14590 38440 -11470
rect 39160 -14590 39200 -11470
rect 38400 -14630 39200 -14590
rect 40000 -11470 40800 -11430
rect 40000 -14590 40040 -11470
rect 40760 -14590 40800 -11470
rect 40000 -14630 40800 -14590
rect 41600 -11470 42400 -11430
rect 41600 -14590 41640 -11470
rect 42360 -14590 42400 -11470
rect 41600 -14630 42400 -14590
rect 43200 -11470 44000 -11430
rect 43200 -14590 43240 -11470
rect 43960 -14590 44000 -11470
rect 43200 -14630 44000 -14590
rect 44800 -11470 45600 -11430
rect 44800 -14590 44840 -11470
rect 45560 -14590 45600 -11470
rect 44800 -14630 45600 -14590
rect 46400 -11470 47200 -11430
rect 46400 -14590 46440 -11470
rect 47160 -14590 47200 -11470
rect 46400 -14630 47200 -14590
<< ndiffc >>
rect -760 50 -40 3170
rect 840 50 1560 3170
rect 2440 50 3160 3170
rect 4040 50 4760 3170
rect 5640 50 6360 3170
rect 7240 50 7960 3170
rect 8840 50 9560 3170
rect 10440 50 11160 3170
rect 12040 50 12760 3170
rect 13640 50 14360 3170
rect 15240 50 15960 3170
rect 16840 50 17560 3170
rect 18440 50 19160 3170
rect 20040 50 20760 3170
rect 21640 50 22360 3170
rect 23240 50 23960 3170
rect 24840 50 25560 3170
rect 26440 50 27160 3170
rect 28040 50 28760 3170
rect 29640 50 30360 3170
rect 31240 50 31960 3170
rect 32840 50 33560 3170
rect 36840 50 37560 3170
rect 38440 50 39160 3170
rect 40040 50 40760 3170
rect 41640 50 42360 3170
rect 43240 50 43960 3170
rect 44840 50 45560 3170
rect 46440 50 47160 3170
rect -760 -4750 -40 -1630
rect 840 -4750 1560 -1630
rect 2440 -4750 3160 -1630
rect 4040 -4750 4760 -1630
rect 5640 -4750 6360 -1630
rect 7240 -4750 7960 -1630
rect 8840 -4750 9560 -1630
rect 10440 -4750 11160 -1630
rect 12040 -4750 12760 -1630
rect 13640 -4750 14360 -1630
rect 15240 -4750 15960 -1630
rect 16840 -4750 17560 -1630
rect 18440 -4750 19160 -1630
rect 20040 -4750 20760 -1630
rect 21640 -4750 22360 -1630
rect 23240 -4750 23960 -1630
rect 24840 -4750 25560 -1630
rect 26440 -4750 27160 -1630
rect 28040 -4750 28760 -1630
rect 29640 -4750 30360 -1630
rect 31240 -4750 31960 -1630
rect 32840 -4750 33560 -1630
rect 36840 -4750 37560 -1630
rect 38440 -4750 39160 -1630
rect 40040 -4750 40760 -1630
rect 41640 -4750 42360 -1630
rect 43240 -4750 43960 -1630
rect 44840 -4750 45560 -1630
rect 46440 -4750 47160 -1630
rect -760 -9790 -40 -6670
rect 840 -9790 1560 -6670
rect 2440 -9790 3160 -6670
rect 4040 -9790 4760 -6670
rect 5640 -9790 6360 -6670
rect 7240 -9790 7960 -6670
rect 8840 -9790 9560 -6670
rect 10440 -9790 11160 -6670
rect 12040 -9790 12760 -6670
rect 13640 -9790 14360 -6670
rect 15240 -9790 15960 -6670
rect 16840 -9790 17560 -6670
rect 18440 -9790 19160 -6670
rect 20040 -9790 20760 -6670
rect 21640 -9790 22360 -6670
rect 23240 -9790 23960 -6670
rect 24840 -9790 25560 -6670
rect 26440 -9790 27160 -6670
rect 28040 -9790 28760 -6670
rect 29640 -9790 30360 -6670
rect 31240 -9790 31960 -6670
rect 32840 -9790 33560 -6670
rect 36840 -9790 37560 -6670
rect 38440 -9790 39160 -6670
rect 40040 -9790 40760 -6670
rect 41640 -9790 42360 -6670
rect 43240 -9790 43960 -6670
rect 44840 -9790 45560 -6670
rect 46440 -9790 47160 -6670
rect -760 -14590 -40 -11470
rect 840 -14590 1560 -11470
rect 2440 -14590 3160 -11470
rect 4040 -14590 4760 -11470
rect 5640 -14590 6360 -11470
rect 7240 -14590 7960 -11470
rect 8840 -14590 9560 -11470
rect 10440 -14590 11160 -11470
rect 12040 -14590 12760 -11470
rect 13640 -14590 14360 -11470
rect 15240 -14590 15960 -11470
rect 16840 -14590 17560 -11470
rect 18440 -14590 19160 -11470
rect 20040 -14590 20760 -11470
rect 21640 -14590 22360 -11470
rect 23240 -14590 23960 -11470
rect 24840 -14590 25560 -11470
rect 26440 -14590 27160 -11470
rect 28040 -14590 28760 -11470
rect 29640 -14590 30360 -11470
rect 31240 -14590 31960 -11470
rect 32840 -14590 33560 -11470
rect 36840 -14590 37560 -11470
rect 38440 -14590 39160 -11470
rect 40040 -14590 40760 -11470
rect 41640 -14590 42360 -11470
rect 43240 -14590 43960 -11470
rect 44840 -14590 45560 -11470
rect 46440 -14590 47160 -11470
<< psubdiff >>
rect -1600 3170 -800 3210
rect -1600 50 -1560 3170
rect -840 50 -800 3170
rect -1600 10 -800 50
rect 22400 3170 23200 3210
rect 22400 50 22440 3170
rect 23160 50 23200 3170
rect 22400 10 23200 50
rect 33600 3170 34400 3210
rect 33600 50 33640 3170
rect 34360 50 34400 3170
rect 33600 10 34400 50
rect 36000 3170 36800 3210
rect 36000 50 36040 3170
rect 36760 50 36800 3170
rect 36000 10 36800 50
rect 47200 3170 48000 3210
rect 47200 50 47240 3170
rect 47960 50 48000 3170
rect 47200 10 48000 50
rect -1600 -1630 -800 -1590
rect -1600 -4750 -1560 -1630
rect -840 -4750 -800 -1630
rect -1600 -4790 -800 -4750
rect 22400 -1630 23200 -1590
rect 22400 -4750 22440 -1630
rect 23160 -4750 23200 -1630
rect 22400 -4790 23200 -4750
rect 33600 -1630 34400 -1590
rect 33600 -4750 33640 -1630
rect 34360 -4750 34400 -1630
rect 33600 -4790 34400 -4750
rect 36000 -1630 36800 -1590
rect 36000 -4750 36040 -1630
rect 36760 -4750 36800 -1630
rect 36000 -4790 36800 -4750
rect 47200 -1630 48000 -1590
rect 47200 -4750 47240 -1630
rect 47960 -4750 48000 -1630
rect 47200 -4790 48000 -4750
rect -1600 -6670 -800 -6630
rect -1600 -9790 -1560 -6670
rect -840 -9790 -800 -6670
rect -1600 -9830 -800 -9790
rect 22400 -6670 23200 -6630
rect 22400 -9790 22440 -6670
rect 23160 -9790 23200 -6670
rect 22400 -9830 23200 -9790
rect 33600 -6670 34400 -6630
rect 33600 -9790 33640 -6670
rect 34360 -9790 34400 -6670
rect 33600 -9830 34400 -9790
rect 36000 -6670 36800 -6630
rect 36000 -9790 36040 -6670
rect 36760 -9790 36800 -6670
rect 36000 -9830 36800 -9790
rect 47200 -6670 48000 -6630
rect 47200 -9790 47240 -6670
rect 47960 -9790 48000 -6670
rect 47200 -9830 48000 -9790
rect -1600 -11470 -800 -11430
rect -1600 -14590 -1560 -11470
rect -840 -14590 -800 -11470
rect -1600 -14630 -800 -14590
rect 22400 -11470 23200 -11430
rect 22400 -14590 22440 -11470
rect 23160 -14590 23200 -11470
rect 22400 -14630 23200 -14590
rect 33600 -11470 34400 -11430
rect 33600 -14590 33640 -11470
rect 34360 -14590 34400 -11470
rect 33600 -14630 34400 -14590
rect 36000 -11470 36800 -11430
rect 36000 -14590 36040 -11470
rect 36760 -14590 36800 -11470
rect 36000 -14630 36800 -14590
rect 47200 -11470 48000 -11430
rect 47200 -14590 47240 -11470
rect 47960 -14590 48000 -11470
rect 47200 -14630 48000 -14590
<< psubdiffcont >>
rect -1560 50 -840 3170
rect 22440 50 23160 3170
rect 33640 50 34360 3170
rect 36040 50 36760 3170
rect 47240 50 47960 3170
rect -1560 -4750 -840 -1630
rect 22440 -4750 23160 -1630
rect 33640 -4750 34360 -1630
rect 36040 -4750 36760 -1630
rect 47240 -4750 47960 -1630
rect -1560 -9790 -840 -6670
rect 22440 -9790 23160 -6670
rect 33640 -9790 34360 -6670
rect 36040 -9790 36760 -6670
rect 47240 -9790 47960 -6670
rect -1560 -14590 -840 -11470
rect 22440 -14590 23160 -11470
rect 33640 -14590 34360 -11470
rect 36040 -14590 36760 -11470
rect 47240 -14590 47960 -11470
<< poly >>
rect 6400 3420 7200 3440
rect 6400 3260 6440 3420
rect 7160 3260 7200 3420
rect 0 3210 800 3240
rect 1600 3210 2400 3240
rect 3200 3210 4000 3240
rect 4800 3210 5600 3240
rect 6400 3210 7200 3260
rect 14400 3420 15200 3440
rect 14400 3260 14440 3420
rect 15160 3260 15200 3420
rect 8000 3210 8800 3240
rect 9600 3210 10400 3240
rect 11200 3210 12000 3240
rect 12800 3210 13600 3240
rect 14400 3210 15200 3260
rect 16000 3210 16800 3240
rect 17600 3210 18400 3240
rect 19200 3210 20000 3240
rect 20800 3210 21600 3240
rect 24000 3210 24800 3240
rect 25600 3210 26400 3240
rect 27200 3210 28000 3240
rect 28800 3210 29600 3240
rect 30400 3210 31200 3240
rect 32000 3210 32800 3240
rect 37600 3210 38400 3240
rect 39200 3210 40000 3240
rect 40800 3210 41600 3240
rect 42400 3210 43200 3240
rect 44000 3210 44800 3240
rect 45600 3210 46400 3240
rect 0 -20 800 10
rect 1600 -20 2400 10
rect 3200 -20 4000 10
rect 4800 -20 5600 10
rect 6400 -20 7200 10
rect 8000 -20 8800 10
rect 9600 -20 10400 10
rect 11200 -20 12000 10
rect 12800 -20 13600 10
rect 14400 -20 15200 10
rect 16000 -20 16800 10
rect 17600 -20 18400 10
rect 19200 -20 20000 10
rect 20800 -20 21600 10
rect 24000 -20 24800 10
rect -780 -40 2400 -20
rect -780 -200 -760 -40
rect -40 -200 840 -40
rect 1560 -200 2400 -40
rect -780 -220 2400 -200
rect 19200 -40 22380 -20
rect 19200 -200 20040 -40
rect 20760 -200 21640 -40
rect 22360 -200 22380 -40
rect 19200 -220 22380 -200
rect 23220 -40 24800 -20
rect 23220 -200 23240 -40
rect 23960 -200 24800 -40
rect 23220 -220 24800 -200
rect 6400 -1380 7200 -1360
rect 6400 -1540 6440 -1380
rect 7160 -1540 7200 -1380
rect 0 -1590 800 -1560
rect 1600 -1590 2400 -1560
rect 3200 -1590 4000 -1560
rect 4800 -1590 5600 -1560
rect 6400 -1590 7200 -1540
rect 14400 -1380 15200 -1360
rect 14400 -1540 14440 -1380
rect 15160 -1540 15200 -1380
rect 8000 -1590 8800 -1560
rect 9600 -1590 10400 -1560
rect 11200 -1590 12000 -1560
rect 12800 -1590 13600 -1560
rect 14400 -1590 15200 -1540
rect 16000 -1590 16800 -1560
rect 17600 -1590 18400 -1560
rect 19200 -1590 20000 -1560
rect 20800 -1590 21600 -1560
rect 24000 -1590 24800 -1560
rect 25600 -1590 26400 10
rect 27200 -1590 28000 10
rect 28800 -1590 29600 10
rect 30400 -1590 31200 10
rect 32000 -20 32800 10
rect 37600 -20 38400 10
rect 32000 -40 33580 -20
rect 32000 -200 32840 -40
rect 33560 -200 33580 -40
rect 32000 -220 33580 -200
rect 36820 -40 38400 -20
rect 36820 -200 36840 -40
rect 37560 -200 38400 -40
rect 36820 -220 38400 -200
rect 32000 -1590 32800 -1560
rect 37600 -1590 38400 -1560
rect 39200 -1590 40000 10
rect 40800 -1590 41600 10
rect 42400 -1590 43200 10
rect 44000 -1590 44800 10
rect 45600 -20 46400 10
rect 45600 -40 47180 -20
rect 45600 -200 46440 -40
rect 47160 -200 47180 -40
rect 45600 -220 47180 -200
rect 45600 -1590 46400 -1560
rect 0 -4820 800 -4790
rect 1600 -4820 2400 -4790
rect 3200 -4820 4000 -4790
rect 4800 -4820 5600 -4790
rect 6400 -4820 7200 -4790
rect 8000 -4820 8800 -4790
rect 9600 -4820 10400 -4790
rect 11200 -4820 12000 -4790
rect 12800 -4820 13600 -4790
rect 14400 -4820 15200 -4790
rect 16000 -4820 16800 -4790
rect 17600 -4820 18400 -4790
rect 19200 -4820 20000 -4790
rect 20800 -4820 21600 -4790
rect 24000 -4820 24800 -4790
rect 25600 -4820 26400 -4790
rect 27200 -4820 28000 -4790
rect 28800 -4820 29600 -4790
rect 30400 -4820 31200 -4790
rect 32000 -4820 32800 -4790
rect 37600 -4820 38400 -4790
rect -780 -4840 2400 -4820
rect -780 -5000 -760 -4840
rect -40 -5000 840 -4840
rect 1560 -5000 2400 -4840
rect -780 -5020 2400 -5000
rect 19200 -4840 22380 -4820
rect 19200 -5000 20040 -4840
rect 20760 -5000 21640 -4840
rect 22360 -5000 22380 -4840
rect 19200 -5020 22380 -5000
rect 23220 -4840 24800 -4820
rect 23220 -5000 23240 -4840
rect 23960 -5000 24800 -4840
rect 23220 -5020 24800 -5000
rect 32000 -4840 33580 -4820
rect 32000 -5000 32840 -4840
rect 33560 -5000 33580 -4840
rect 32000 -5020 33580 -5000
rect 36820 -4840 38400 -4820
rect 36820 -5000 36840 -4840
rect 37560 -5000 38400 -4840
rect 36820 -5020 38400 -5000
rect 0 -6630 800 -6600
rect 1600 -6630 2400 -6600
rect 3200 -6630 4000 -6600
rect 4800 -6630 5600 -6600
rect 6400 -6630 7200 -6600
rect 8000 -6630 8800 -6600
rect 9600 -6630 10400 -6600
rect 11200 -6630 12000 -6600
rect 12800 -6630 13600 -6600
rect 14400 -6630 15200 -6600
rect 16000 -6630 16800 -6600
rect 17600 -6630 18400 -6600
rect 19200 -6630 20000 -6600
rect 20800 -6630 21600 -6600
rect 24000 -6630 24800 -6600
rect 25600 -6630 26400 -6600
rect 27200 -6630 28000 -6600
rect 28800 -6630 29600 -6600
rect 30400 -6630 31200 -6600
rect 32000 -6630 32800 -6600
rect 37600 -6630 38400 -6600
rect 39200 -6630 40000 -4790
rect 40800 -6630 41600 -4790
rect 42400 -6630 43200 -4790
rect 44000 -6630 44800 -4790
rect 45600 -4820 46400 -4790
rect 45600 -4840 47180 -4820
rect 45600 -5000 46440 -4840
rect 47160 -5000 47180 -4840
rect 45600 -5020 47180 -5000
rect 45600 -6630 46400 -6600
rect 0 -9860 800 -9830
rect -780 -9880 800 -9860
rect -780 -10040 -760 -9880
rect -40 -10040 800 -9880
rect -780 -10060 800 -10040
rect 1600 -9860 2400 -9830
rect 3200 -9860 4000 -9830
rect 4800 -9860 5600 -9830
rect 6400 -9860 7200 -9830
rect 8000 -9860 8800 -9830
rect 9600 -9860 10400 -9830
rect 11200 -9860 12000 -9830
rect 12800 -9860 13600 -9830
rect 14400 -9860 15200 -9830
rect 16000 -9860 16800 -9830
rect 17600 -9860 18400 -9830
rect 19200 -9860 20000 -9830
rect 20800 -9860 21600 -9830
rect 24000 -9860 24800 -9830
rect 1600 -11240 1630 -9860
rect 3200 -11240 3230 -9860
rect 4800 -11240 4830 -9860
rect 6400 -11240 6430 -9860
rect 8000 -9880 8900 -9860
rect 8000 -9920 8840 -9880
rect 8880 -9920 8900 -9880
rect 8000 -9940 8900 -9920
rect 9600 -11240 9630 -9860
rect 11200 -11240 11230 -9860
rect 13170 -9880 13250 -9860
rect 13170 -9920 13190 -9880
rect 13230 -9920 13250 -9880
rect 13170 -9940 13250 -9920
rect 14400 -11240 14430 -9860
rect 16000 -11240 16030 -9860
rect 17600 -11240 17630 -9860
rect 19200 -11240 19230 -9860
rect 20800 -9880 22380 -9860
rect 20800 -10040 21640 -9880
rect 22360 -10040 22380 -9880
rect 20800 -10060 22380 -10040
rect 23220 -9880 24800 -9860
rect 23220 -10040 23240 -9880
rect 23960 -10040 24800 -9880
rect 23220 -10060 24800 -10040
rect 1600 -11270 12000 -11240
rect 1600 -11290 2500 -11270
rect 1600 -11330 2440 -11290
rect 2480 -11330 2500 -11290
rect 1600 -11350 2500 -11330
rect 3200 -11290 4100 -11270
rect 3200 -11330 4040 -11290
rect 4080 -11330 4100 -11290
rect 3200 -11350 4100 -11330
rect 4800 -11290 5700 -11270
rect 4800 -11330 5640 -11290
rect 5680 -11330 5700 -11290
rect 4800 -11350 5700 -11330
rect 0 -11430 800 -11400
rect 1600 -11430 2400 -11350
rect 3200 -11430 4000 -11350
rect 4800 -11430 5600 -11350
rect 6400 -11430 7200 -11270
rect 8000 -11340 8900 -11320
rect 8000 -11380 8840 -11340
rect 8880 -11380 8900 -11340
rect 8000 -11400 8900 -11380
rect 8000 -11430 8800 -11400
rect 9600 -11430 10400 -11270
rect 11200 -11430 12000 -11270
rect 14400 -11270 23200 -11240
rect 13170 -11340 13250 -11320
rect 13170 -11380 13190 -11340
rect 13230 -11380 13250 -11340
rect 13170 -11400 13250 -11380
rect 12800 -11430 13600 -11400
rect 14400 -11430 15200 -11270
rect 16000 -11430 16800 -11270
rect 17600 -11430 18400 -11270
rect 19200 -11290 20100 -11270
rect 19200 -11330 20040 -11290
rect 20080 -11330 20100 -11290
rect 19200 -11350 20100 -11330
rect 19200 -11430 20000 -11350
rect 20800 -11430 21600 -11400
rect 24000 -11430 24800 -11400
rect 25600 -11430 26400 -9830
rect 27200 -11430 28000 -9830
rect 28800 -11430 29600 -9830
rect 30400 -11430 31200 -9830
rect 32000 -9860 32800 -9830
rect 37600 -9860 38400 -9830
rect 39200 -9860 40000 -9830
rect 40800 -9860 41600 -9830
rect 42400 -9860 43200 -9830
rect 44000 -9860 44800 -9830
rect 45600 -9860 46400 -9830
rect 32000 -9880 33580 -9860
rect 32000 -10040 32840 -9880
rect 33560 -10040 33580 -9880
rect 32000 -10060 33580 -10040
rect 36820 -9880 38400 -9860
rect 36820 -10040 36840 -9880
rect 37560 -10040 38400 -9880
rect 36820 -10060 38400 -10040
rect 45600 -9880 47180 -9860
rect 45600 -10040 46440 -9880
rect 47160 -10040 47180 -9880
rect 45600 -10060 47180 -10040
rect 32000 -11430 32800 -11400
rect 37600 -11430 38400 -11400
rect 39200 -11430 40000 -11400
rect 40800 -11430 41600 -11400
rect 42400 -11430 43200 -11400
rect 44000 -11430 44800 -11400
rect 45600 -11430 46400 -11400
rect 0 -14660 800 -14630
rect 1600 -14660 2400 -14630
rect 3200 -14660 4000 -14630
rect 4800 -14660 5600 -14630
rect 6400 -14660 7200 -14630
rect 8000 -14660 8800 -14630
rect 9600 -14660 10400 -14630
rect 11200 -14660 12000 -14630
rect 12800 -14660 13600 -14630
rect -780 -14680 800 -14660
rect -780 -14840 -760 -14680
rect -40 -14840 800 -14680
rect -780 -14860 800 -14840
rect 14400 -14680 15200 -14630
rect 14400 -14840 14420 -14680
rect 15180 -14840 15200 -14680
rect 14400 -14860 15200 -14840
rect 16000 -14680 16800 -14630
rect 16000 -14840 16020 -14680
rect 16780 -14840 16800 -14680
rect 16000 -14860 16800 -14840
rect 17600 -14680 18400 -14630
rect 17600 -14840 17620 -14680
rect 18380 -14840 18400 -14680
rect 17600 -14860 18400 -14840
rect 19200 -14680 20000 -14630
rect 19200 -14840 19220 -14680
rect 19980 -14840 20000 -14680
rect 19200 -14860 20000 -14840
rect 20800 -14660 21600 -14630
rect 24000 -14660 24800 -14630
rect 20800 -14680 22380 -14660
rect 20800 -14840 21640 -14680
rect 22360 -14840 22380 -14680
rect 20800 -14860 22380 -14840
rect 23220 -14680 24800 -14660
rect 23220 -14840 23240 -14680
rect 23960 -14840 24800 -14680
rect 23220 -14860 24800 -14840
rect 25600 -14680 26400 -14630
rect 25600 -14840 25620 -14680
rect 26380 -14840 26400 -14680
rect 25600 -14860 26400 -14840
rect 27200 -14680 28000 -14630
rect 28800 -14660 29600 -14630
rect 30400 -14660 31200 -14630
rect 32000 -14660 32800 -14630
rect 37600 -14660 38400 -14630
rect 27200 -14840 27220 -14680
rect 27980 -14840 28000 -14680
rect 27200 -14860 28000 -14840
rect 32000 -14680 33580 -14660
rect 32000 -14840 32840 -14680
rect 33560 -14840 33580 -14680
rect 32000 -14860 33580 -14840
rect 36820 -14680 38400 -14660
rect 36820 -14840 36840 -14680
rect 37560 -14840 38400 -14680
rect 36820 -14860 38400 -14840
rect 39200 -14680 40000 -14630
rect 39200 -14840 39220 -14680
rect 39980 -14840 40000 -14680
rect 39200 -14860 40000 -14840
rect 40800 -14680 41600 -14630
rect 40800 -14840 40820 -14680
rect 41580 -14840 41600 -14680
rect 40800 -14860 41600 -14840
rect 42400 -14680 43200 -14630
rect 42400 -14840 42420 -14680
rect 43180 -14840 43200 -14680
rect 42400 -14860 43200 -14840
rect 44000 -14680 44800 -14630
rect 44000 -14840 44020 -14680
rect 44780 -14840 44800 -14680
rect 44000 -14860 44800 -14840
rect 45600 -14660 46400 -14630
rect 45600 -14680 47180 -14660
rect 45600 -14840 46440 -14680
rect 47160 -14840 47180 -14680
rect 45600 -14860 47180 -14840
<< polycont >>
rect 6440 3260 7160 3420
rect 14440 3260 15160 3420
rect -760 -200 -40 -40
rect 840 -200 1560 -40
rect 20040 -200 20760 -40
rect 21640 -200 22360 -40
rect 23240 -200 23960 -40
rect 6440 -1540 7160 -1380
rect 14440 -1540 15160 -1380
rect 32840 -200 33560 -40
rect 36840 -200 37560 -40
rect 46440 -200 47160 -40
rect -760 -5000 -40 -4840
rect 840 -5000 1560 -4840
rect 20040 -5000 20760 -4840
rect 21640 -5000 22360 -4840
rect 23240 -5000 23960 -4840
rect 32840 -5000 33560 -4840
rect 36840 -5000 37560 -4840
rect 46440 -5000 47160 -4840
rect -760 -10040 -40 -9880
rect 8840 -9920 8880 -9880
rect 13190 -9920 13230 -9880
rect 21640 -10040 22360 -9880
rect 23240 -10040 23960 -9880
rect 2440 -11330 2480 -11290
rect 4040 -11330 4080 -11290
rect 5640 -11330 5680 -11290
rect 8840 -11380 8880 -11340
rect 13190 -11380 13230 -11340
rect 20040 -11330 20080 -11290
rect 32840 -10040 33560 -9880
rect 36840 -10040 37560 -9880
rect 46440 -10040 47160 -9880
rect -760 -14840 -40 -14680
rect 14420 -14840 15180 -14680
rect 16020 -14840 16780 -14680
rect 17620 -14840 18380 -14680
rect 19220 -14840 19980 -14680
rect 21640 -14840 22360 -14680
rect 23240 -14840 23960 -14680
rect 25620 -14840 26380 -14680
rect 27220 -14840 27980 -14680
rect 32840 -14840 33560 -14680
rect 36840 -14840 37560 -14680
rect 39220 -14840 39980 -14680
rect 40820 -14840 41580 -14680
rect 42420 -14840 43180 -14680
rect 44020 -14840 44780 -14680
rect 46440 -14840 47160 -14680
<< locali >>
rect 6420 3420 7180 3440
rect 6420 3260 6440 3420
rect 7160 3260 7180 3420
rect 6420 3240 7180 3260
rect 14420 3420 15180 3440
rect 14420 3260 14440 3420
rect 15160 3260 15180 3420
rect 14420 3240 15180 3260
rect 40400 3290 43600 3490
rect 40400 3190 40780 3290
rect 43220 3190 43600 3290
rect -1580 3170 -20 3190
rect -1580 50 -1560 3170
rect -840 50 -760 3170
rect -40 50 -20 3170
rect -1580 30 -20 50
rect -780 -40 -20 30
rect -780 -200 -760 -40
rect -40 -200 -20 -40
rect -780 -220 -20 -200
rect 820 3170 1580 3190
rect 820 50 840 3170
rect 1560 50 1580 3170
rect 820 -40 1580 50
rect 2420 3170 3180 3190
rect 2420 50 2440 3170
rect 3160 50 3180 3170
rect 2420 30 3180 50
rect 4020 3170 4780 3190
rect 4020 50 4040 3170
rect 4760 50 4780 3170
rect 4020 30 4780 50
rect 5620 3170 6380 3190
rect 5620 50 5640 3170
rect 6360 50 6380 3170
rect 5620 30 6380 50
rect 7220 3170 7980 3190
rect 7220 50 7240 3170
rect 7960 50 7980 3170
rect 7220 30 7980 50
rect 8820 3170 9580 3190
rect 8820 50 8840 3170
rect 9560 50 9580 3170
rect 8820 30 9580 50
rect 10420 3170 11180 3190
rect 10420 50 10440 3170
rect 11160 50 11180 3170
rect 10420 30 11180 50
rect 12020 3170 12780 3190
rect 12020 50 12040 3170
rect 12760 50 12780 3170
rect 12020 30 12780 50
rect 13620 3170 14380 3190
rect 13620 50 13640 3170
rect 14360 50 14380 3170
rect 13620 30 14380 50
rect 15220 3170 15980 3190
rect 15220 50 15240 3170
rect 15960 50 15980 3170
rect 15220 30 15980 50
rect 16820 3170 17580 3190
rect 16820 50 16840 3170
rect 17560 50 17580 3170
rect 16820 30 17580 50
rect 18420 3170 19180 3190
rect 18420 50 18440 3170
rect 19160 50 19180 3170
rect 18420 30 19180 50
rect 20020 3170 20780 3190
rect 20020 50 20040 3170
rect 20760 50 20780 3170
rect 820 -200 840 -40
rect 1560 -200 1580 -40
rect 820 -220 1580 -200
rect 20020 -40 20780 50
rect 20020 -200 20040 -40
rect 20760 -200 20780 -40
rect 20020 -220 20780 -200
rect 21620 3170 23980 3190
rect 21620 50 21640 3170
rect 22360 50 22440 3170
rect 23160 50 23240 3170
rect 23960 50 23980 3170
rect 21620 30 23980 50
rect 24820 3170 25580 3190
rect 24820 50 24840 3170
rect 25560 50 25580 3170
rect 24820 30 25580 50
rect 26420 3170 27180 3190
rect 26420 50 26440 3170
rect 27160 50 27180 3170
rect 26420 30 27180 50
rect 28020 3170 28780 3190
rect 28020 50 28040 3170
rect 28760 50 28780 3170
rect 28020 30 28780 50
rect 29620 3170 30380 3190
rect 29620 50 29640 3170
rect 30360 50 30380 3170
rect 29620 30 30380 50
rect 31220 3170 31980 3190
rect 31220 50 31240 3170
rect 31960 50 31980 3170
rect 31220 30 31980 50
rect 32820 3170 34380 3190
rect 32820 50 32840 3170
rect 33560 50 33640 3170
rect 34360 50 34380 3170
rect 32820 30 34380 50
rect 36020 3170 37580 3190
rect 36020 50 36040 3170
rect 36760 50 36840 3170
rect 37560 50 37580 3170
rect 36020 30 37580 50
rect 38420 3170 39180 3190
rect 38420 50 38440 3170
rect 39160 50 39180 3170
rect 38420 30 39180 50
rect 40020 3170 40780 3190
rect 40020 50 40040 3170
rect 40760 50 40780 3170
rect 40020 30 40780 50
rect 41620 3170 42380 3190
rect 41620 50 41640 3170
rect 42360 50 42380 3170
rect 41620 30 42380 50
rect 43220 3170 43980 3190
rect 43220 50 43240 3170
rect 43960 50 43980 3170
rect 43220 30 43980 50
rect 44820 3170 45580 3190
rect 44820 50 44840 3170
rect 45560 50 45580 3170
rect 44820 30 45580 50
rect 46420 3170 47980 3190
rect 46420 50 46440 3170
rect 47160 50 47240 3170
rect 47960 50 47980 3170
rect 46420 30 47980 50
rect 21620 -40 22380 30
rect 21620 -200 21640 -40
rect 22360 -200 22380 -40
rect 21620 -220 22380 -200
rect 23220 -40 23980 30
rect 23220 -200 23240 -40
rect 23960 -200 23980 -40
rect 23220 -220 23980 -200
rect 32820 -40 33580 30
rect 32820 -200 32840 -40
rect 33560 -200 33580 -40
rect 32820 -220 33580 -200
rect 36820 -40 37580 30
rect 36820 -200 36840 -40
rect 37560 -200 37580 -40
rect 36820 -220 37580 -200
rect 46420 -40 47180 30
rect 46420 -200 46440 -40
rect 47160 -200 47180 -40
rect 46420 -220 47180 -200
rect 6420 -1380 7180 -1360
rect 6420 -1540 6440 -1380
rect 7160 -1540 7180 -1380
rect 6420 -1560 7180 -1540
rect 14420 -1380 15180 -1360
rect 14420 -1540 14440 -1380
rect 15160 -1540 15180 -1380
rect 14420 -1560 15180 -1540
rect 40400 -1510 43600 -1310
rect 40400 -1610 40780 -1510
rect 43220 -1610 43600 -1510
rect -1580 -1630 -20 -1610
rect -1580 -4750 -1560 -1630
rect -840 -4750 -760 -1630
rect -40 -4750 -20 -1630
rect -1580 -4770 -20 -4750
rect -780 -4840 -20 -4770
rect -780 -5000 -760 -4840
rect -40 -5000 -20 -4840
rect -780 -5020 -20 -5000
rect 820 -1630 1580 -1610
rect 820 -4750 840 -1630
rect 1560 -4750 1580 -1630
rect 820 -4840 1580 -4750
rect 2420 -1630 3180 -1610
rect 2420 -4750 2440 -1630
rect 3160 -4750 3180 -1630
rect 2420 -4770 3180 -4750
rect 4020 -1630 4780 -1610
rect 4020 -4750 4040 -1630
rect 4760 -4750 4780 -1630
rect 4020 -4770 4780 -4750
rect 5620 -1630 6380 -1610
rect 5620 -4750 5640 -1630
rect 6360 -4750 6380 -1630
rect 5620 -4770 6380 -4750
rect 7220 -1630 7980 -1610
rect 7220 -4750 7240 -1630
rect 7960 -4750 7980 -1630
rect 7220 -4770 7980 -4750
rect 8820 -1630 9580 -1610
rect 8820 -4750 8840 -1630
rect 9560 -4750 9580 -1630
rect 8820 -4770 9580 -4750
rect 10420 -1630 11180 -1610
rect 10420 -4750 10440 -1630
rect 11160 -4750 11180 -1630
rect 10420 -4770 11180 -4750
rect 12020 -1630 12780 -1610
rect 12020 -4750 12040 -1630
rect 12760 -4750 12780 -1630
rect 12020 -4770 12780 -4750
rect 13620 -1630 14380 -1610
rect 13620 -4750 13640 -1630
rect 14360 -4750 14380 -1630
rect 13620 -4770 14380 -4750
rect 15220 -1630 15980 -1610
rect 15220 -4750 15240 -1630
rect 15960 -4750 15980 -1630
rect 15220 -4770 15980 -4750
rect 16820 -1630 17580 -1610
rect 16820 -4750 16840 -1630
rect 17560 -4750 17580 -1630
rect 16820 -4770 17580 -4750
rect 18420 -1630 19180 -1610
rect 18420 -4750 18440 -1630
rect 19160 -4750 19180 -1630
rect 18420 -4770 19180 -4750
rect 20020 -1630 20780 -1610
rect 20020 -4750 20040 -1630
rect 20760 -4750 20780 -1630
rect 820 -5000 840 -4840
rect 1560 -5000 1580 -4840
rect 820 -5020 1580 -5000
rect 20020 -4840 20780 -4750
rect 20020 -5000 20040 -4840
rect 20760 -5000 20780 -4840
rect 20020 -5020 20780 -5000
rect 21620 -1630 23980 -1610
rect 21620 -4750 21640 -1630
rect 22360 -4750 22440 -1630
rect 23160 -4750 23240 -1630
rect 23960 -4750 23980 -1630
rect 21620 -4770 23980 -4750
rect 24820 -1630 25580 -1610
rect 24820 -4750 24840 -1630
rect 25560 -4750 25580 -1630
rect 24820 -4770 25580 -4750
rect 26420 -1630 27180 -1610
rect 26420 -4750 26440 -1630
rect 27160 -4750 27180 -1630
rect 26420 -4770 27180 -4750
rect 28020 -1630 28780 -1610
rect 28020 -4750 28040 -1630
rect 28760 -4750 28780 -1630
rect 28020 -4770 28780 -4750
rect 29620 -1630 30380 -1610
rect 29620 -4750 29640 -1630
rect 30360 -4750 30380 -1630
rect 29620 -4770 30380 -4750
rect 31220 -1630 31980 -1610
rect 31220 -4750 31240 -1630
rect 31960 -4750 31980 -1630
rect 31220 -4770 31980 -4750
rect 32820 -1630 34380 -1610
rect 32820 -4750 32840 -1630
rect 33560 -4750 33640 -1630
rect 34360 -4750 34380 -1630
rect 32820 -4770 34380 -4750
rect 36020 -1630 37580 -1610
rect 36020 -4750 36040 -1630
rect 36760 -4750 36840 -1630
rect 37560 -4750 37580 -1630
rect 36020 -4770 37580 -4750
rect 38420 -1630 39180 -1610
rect 38420 -4750 38440 -1630
rect 39160 -4750 39180 -1630
rect 38420 -4770 39180 -4750
rect 40020 -1630 40780 -1610
rect 40020 -4750 40040 -1630
rect 40760 -4750 40780 -1630
rect 40020 -4770 40780 -4750
rect 41620 -1630 42380 -1610
rect 41620 -4750 41640 -1630
rect 42360 -4750 42380 -1630
rect 41620 -4770 42380 -4750
rect 43220 -1630 43980 -1610
rect 43220 -4750 43240 -1630
rect 43960 -4750 43980 -1630
rect 43220 -4770 43980 -4750
rect 44820 -1630 45580 -1610
rect 44820 -4750 44840 -1630
rect 45560 -4750 45580 -1630
rect 44820 -4770 45580 -4750
rect 46420 -1630 47980 -1610
rect 46420 -4750 46440 -1630
rect 47160 -4750 47240 -1630
rect 47960 -4750 47980 -1630
rect 46420 -4770 47980 -4750
rect 21620 -4840 22380 -4770
rect 21620 -5000 21640 -4840
rect 22360 -5000 22380 -4840
rect 21620 -5020 22380 -5000
rect 23220 -4840 23980 -4770
rect 23220 -5000 23240 -4840
rect 23960 -5000 23980 -4840
rect 23220 -5020 23980 -5000
rect 32820 -4840 33580 -4770
rect 32820 -5000 32840 -4840
rect 33560 -5000 33580 -4840
rect 32820 -5020 33580 -5000
rect 36820 -4840 37580 -4770
rect 36820 -5000 36840 -4840
rect 37560 -5000 37580 -4840
rect 36820 -5020 37580 -5000
rect 46420 -4840 47180 -4770
rect 46420 -5000 46440 -4840
rect 47160 -5000 47180 -4840
rect 46420 -5020 47180 -5000
rect 40400 -6550 43600 -6350
rect 40400 -6650 40780 -6550
rect 43220 -6650 43600 -6550
rect -1580 -6670 -20 -6650
rect -1580 -9790 -1560 -6670
rect -840 -9790 -760 -6670
rect -40 -9790 -20 -6670
rect -1580 -9810 -20 -9790
rect -780 -9880 -20 -9810
rect -780 -10040 -760 -9880
rect -40 -10040 -20 -9880
rect -780 -10060 -20 -10040
rect 820 -6670 1580 -6650
rect 820 -9790 840 -6670
rect 1560 -9790 1580 -6670
rect 820 -9810 1580 -9790
rect 2420 -6670 3180 -6650
rect 2420 -9790 2440 -6670
rect 3160 -9790 3180 -6670
rect 2420 -9810 3180 -9790
rect 4020 -6670 4780 -6650
rect 4020 -9790 4040 -6670
rect 4760 -9790 4780 -6670
rect 4020 -9810 4780 -9790
rect 5620 -6670 6380 -6650
rect 5620 -9790 5640 -6670
rect 6360 -9790 6380 -6670
rect 5620 -9810 6380 -9790
rect 7220 -6670 7980 -6650
rect 7220 -9790 7240 -6670
rect 7960 -9790 7980 -6670
rect 7220 -9810 7980 -9790
rect 8820 -6670 9580 -6650
rect 8820 -9790 8840 -6670
rect 9560 -9790 9580 -6670
rect 820 -10110 860 -9810
rect 4020 -10110 4060 -9810
rect 7220 -10110 7260 -9810
rect 8820 -9860 9580 -9790
rect 10420 -6670 11180 -6650
rect 10420 -9790 10440 -6670
rect 11160 -9790 11180 -6670
rect 10420 -9810 11180 -9790
rect 12020 -6670 12780 -6650
rect 12020 -9790 12040 -6670
rect 12760 -9790 12780 -6670
rect 12020 -9810 12780 -9790
rect 13620 -6670 14380 -6650
rect 13620 -9790 13640 -6670
rect 14360 -9790 14380 -6670
rect 13620 -9810 14380 -9790
rect 15220 -6670 15980 -6650
rect 15220 -9790 15240 -6670
rect 15960 -9790 15980 -6670
rect 15220 -9810 15980 -9790
rect 16820 -6670 17580 -6650
rect 16820 -9790 16840 -6670
rect 17560 -9790 17580 -6670
rect 16820 -9810 17580 -9790
rect 18420 -6670 19180 -6650
rect 18420 -9790 18440 -6670
rect 19160 -9790 19180 -6670
rect 18420 -9810 19180 -9790
rect 20020 -6670 20780 -6650
rect 20020 -9790 20040 -6670
rect 20760 -9790 20780 -6670
rect 20020 -9810 20780 -9790
rect 8820 -9880 8900 -9860
rect 8820 -9920 8840 -9880
rect 8880 -9920 8900 -9880
rect 8820 -9940 8900 -9920
rect -1600 -10150 7260 -10110
rect 820 -11450 860 -10150
rect 2420 -11290 2500 -11270
rect 2420 -11330 2440 -11290
rect 2480 -11330 2500 -11290
rect 2420 -11350 2500 -11330
rect 4020 -11290 4100 -11270
rect 4020 -11330 4040 -11290
rect 4080 -11330 4100 -11290
rect 4020 -11350 4100 -11330
rect 5620 -11290 5700 -11270
rect 5620 -11330 5640 -11290
rect 5680 -11330 5700 -11290
rect 5620 -11350 5700 -11330
rect -1580 -11470 -20 -11450
rect -1580 -14590 -1560 -11470
rect -840 -14590 -760 -11470
rect -40 -14590 -20 -11470
rect -1580 -14610 -20 -14590
rect 820 -11470 1580 -11450
rect 820 -14590 840 -11470
rect 1560 -14590 1580 -11470
rect 820 -14610 1580 -14590
rect 2420 -11470 3180 -11350
rect 2420 -14590 2440 -11470
rect 3160 -14590 3180 -11470
rect 2420 -14610 3180 -14590
rect 4020 -11470 4780 -11350
rect 4020 -14590 4040 -11470
rect 4760 -14590 4780 -11470
rect 4020 -14610 4780 -14590
rect 5620 -11470 6380 -11350
rect 5620 -14590 5640 -11470
rect 6360 -14590 6380 -11470
rect 5620 -14610 6380 -14590
rect 7220 -11450 7260 -10150
rect 8820 -11340 8900 -11320
rect 8820 -11380 8840 -11340
rect 8880 -11380 8900 -11340
rect 8820 -11400 8900 -11380
rect 7220 -11470 7980 -11450
rect 7220 -14590 7240 -11470
rect 7960 -14590 7980 -11470
rect 7220 -14610 7980 -14590
rect 8820 -11470 9580 -11400
rect 8820 -14590 8840 -11470
rect 9560 -14590 9580 -11470
rect 8820 -14610 9580 -14590
rect 10420 -11450 10460 -9810
rect 12020 -11450 12060 -9810
rect 13170 -9880 13330 -9860
rect 13170 -9920 13190 -9880
rect 13230 -9920 13270 -9880
rect 13310 -9920 13330 -9880
rect 13170 -9940 13330 -9920
rect 13170 -11340 13330 -11320
rect 13170 -11380 13190 -11340
rect 13230 -11380 13270 -11340
rect 13310 -11380 13330 -11340
rect 13170 -11400 13330 -11380
rect 13620 -11450 13660 -9810
rect 15220 -11450 15260 -9810
rect 18420 -11450 18460 -9810
rect 20020 -11290 20100 -11270
rect 20020 -11330 20040 -11290
rect 20080 -11330 20100 -11290
rect 20020 -11350 20100 -11330
rect 20740 -11350 20780 -9810
rect 21620 -6670 23980 -6650
rect 21620 -9790 21640 -6670
rect 22360 -9790 22440 -6670
rect 23160 -9790 23240 -6670
rect 23960 -9790 23980 -6670
rect 21620 -9810 23980 -9790
rect 24820 -6670 25580 -6650
rect 24820 -9790 24840 -6670
rect 25560 -9790 25580 -6670
rect 24820 -9810 25580 -9790
rect 26420 -6670 27180 -6650
rect 26420 -9790 26440 -6670
rect 27160 -9790 27180 -6670
rect 26420 -9810 27180 -9790
rect 28020 -6670 28780 -6650
rect 28020 -9790 28040 -6670
rect 28760 -9790 28780 -6670
rect 28020 -9810 28780 -9790
rect 29620 -6670 30380 -6650
rect 29620 -9790 29640 -6670
rect 30360 -9790 30380 -6670
rect 29620 -9810 30380 -9790
rect 31220 -6670 31980 -6650
rect 31220 -9790 31240 -6670
rect 31960 -9790 31980 -6670
rect 31220 -9810 31980 -9790
rect 32820 -6670 34380 -6650
rect 32820 -9790 32840 -6670
rect 33560 -9790 33640 -6670
rect 34360 -9790 34380 -6670
rect 32820 -9810 34380 -9790
rect 36020 -6670 37580 -6650
rect 36020 -9790 36040 -6670
rect 36760 -9790 36840 -6670
rect 37560 -9790 37580 -6670
rect 36020 -9810 37580 -9790
rect 38420 -6670 39180 -6650
rect 38420 -9790 38440 -6670
rect 39160 -9790 39180 -6670
rect 38420 -9810 39180 -9790
rect 40020 -6670 40780 -6650
rect 40020 -9790 40040 -6670
rect 40760 -9790 40780 -6670
rect 40020 -9810 40780 -9790
rect 41620 -6670 42380 -6650
rect 41620 -9790 41640 -6670
rect 42360 -9790 42380 -6670
rect 41620 -9810 42380 -9790
rect 43220 -6670 43980 -6650
rect 43220 -9790 43240 -6670
rect 43960 -9790 43980 -6670
rect 43220 -9810 43980 -9790
rect 44820 -6670 45580 -6650
rect 44820 -9790 44840 -6670
rect 45560 -9790 45580 -6670
rect 44820 -9810 45580 -9790
rect 46420 -6670 47980 -6650
rect 46420 -9790 46440 -6670
rect 47160 -9790 47240 -6670
rect 47960 -9790 47980 -6670
rect 46420 -9810 47980 -9790
rect 21620 -9880 22380 -9810
rect 21620 -10040 21640 -9880
rect 22360 -10040 22380 -9880
rect 21620 -10060 22380 -10040
rect 23220 -9880 23980 -9810
rect 23220 -10040 23240 -9880
rect 23960 -10040 23980 -9880
rect 23220 -10060 23980 -10040
rect 32820 -9880 33580 -9810
rect 32820 -10040 32840 -9880
rect 33560 -10040 33580 -9880
rect 32820 -10060 33580 -10040
rect 36820 -9880 37580 -9810
rect 36820 -10040 36840 -9880
rect 37560 -10040 37580 -9880
rect 36820 -10060 37580 -10040
rect 46420 -9880 47180 -9810
rect 46420 -10040 46440 -9880
rect 47160 -10040 47180 -9880
rect 46420 -10060 47180 -10040
rect 10420 -11470 11180 -11450
rect 10420 -14590 10440 -11470
rect 11160 -14590 11180 -11470
rect 10420 -14610 11180 -14590
rect 12020 -11470 12780 -11450
rect 12020 -14590 12040 -11470
rect 12760 -14590 12780 -11470
rect 12020 -14610 12780 -14590
rect 13620 -11470 14380 -11450
rect 13620 -14590 13640 -11470
rect 14360 -14590 14380 -11470
rect 13620 -14610 14380 -14590
rect 15220 -11470 15980 -11450
rect 15220 -14590 15240 -11470
rect 15960 -14590 15980 -11470
rect 15220 -14610 15980 -14590
rect 16820 -11470 17580 -11450
rect 16820 -14590 16840 -11470
rect 17560 -14590 17580 -11470
rect 16820 -14610 17580 -14590
rect 18420 -11470 19180 -11450
rect 18420 -14590 18440 -11470
rect 19160 -14590 19180 -11470
rect 18420 -14610 19180 -14590
rect 20020 -11470 20780 -11350
rect 40400 -11350 43600 -11150
rect 40400 -11450 40780 -11350
rect 43220 -11450 43600 -11350
rect 20020 -14590 20040 -11470
rect 20760 -14590 20780 -11470
rect 20020 -14610 20780 -14590
rect 21620 -11470 23980 -11450
rect 21620 -14590 21640 -11470
rect 22360 -14590 22440 -11470
rect 23160 -14590 23240 -11470
rect 23960 -14590 23980 -11470
rect 21620 -14610 23980 -14590
rect 24820 -11470 25580 -11450
rect 24820 -14590 24840 -11470
rect 25560 -14590 25580 -11470
rect 24820 -14610 25580 -14590
rect 26420 -11470 27180 -11450
rect 26420 -14590 26440 -11470
rect 27160 -14590 27180 -11470
rect 26420 -14610 27180 -14590
rect 28020 -11470 28780 -11450
rect 28020 -14590 28040 -11470
rect 28760 -14590 28780 -11470
rect 28020 -14610 28780 -14590
rect 29620 -11470 30380 -11450
rect 29620 -14590 29640 -11470
rect 30360 -14590 30380 -11470
rect 29620 -14610 30380 -14590
rect 31220 -11470 31980 -11450
rect 31220 -14590 31240 -11470
rect 31960 -14590 31980 -11470
rect 31220 -14610 31980 -14590
rect 32820 -11470 34380 -11450
rect 32820 -14590 32840 -11470
rect 33560 -14590 33640 -11470
rect 34360 -14590 34380 -11470
rect 32820 -14610 34380 -14590
rect 36020 -11470 37580 -11450
rect 36020 -14590 36040 -11470
rect 36760 -14590 36840 -11470
rect 37560 -14590 37580 -11470
rect 36020 -14610 37580 -14590
rect 38420 -11470 39180 -11450
rect 38420 -14590 38440 -11470
rect 39160 -14590 39180 -11470
rect 38420 -14610 39180 -14590
rect 40020 -11470 40780 -11450
rect 40020 -14590 40040 -11470
rect 40760 -14590 40780 -11470
rect 40020 -14610 40780 -14590
rect 41620 -11470 42380 -11450
rect 41620 -14590 41640 -11470
rect 42360 -14590 42380 -11470
rect 41620 -14610 42380 -14590
rect 43220 -11470 43980 -11450
rect 43220 -14590 43240 -11470
rect 43960 -14590 43980 -11470
rect 43220 -14610 43980 -14590
rect 44820 -11470 45580 -11450
rect 44820 -14590 44840 -11470
rect 45560 -14590 45580 -11470
rect 44820 -14610 45580 -14590
rect 46420 -11470 47980 -11450
rect 46420 -14590 46440 -11470
rect 47160 -14590 47240 -11470
rect 47960 -14590 47980 -11470
rect 46420 -14610 47980 -14590
rect -780 -14680 -20 -14610
rect -780 -14840 -760 -14680
rect -40 -14840 -20 -14680
rect -780 -14860 -20 -14840
rect 14400 -14680 15200 -14660
rect 14400 -14840 14420 -14680
rect 15180 -14840 15200 -14680
rect 14400 -14910 15200 -14840
rect 16000 -14680 16800 -14660
rect 16000 -14840 16020 -14680
rect 16780 -14840 16800 -14680
rect 16000 -14910 16800 -14840
rect 17600 -14680 18400 -14660
rect 17600 -14840 17620 -14680
rect 18380 -14840 18400 -14680
rect 17600 -14910 18400 -14840
rect 19200 -14680 20000 -14660
rect 19200 -14840 19220 -14680
rect 19980 -14840 20000 -14680
rect 19200 -14910 20000 -14840
rect 21620 -14680 22380 -14610
rect 21620 -14840 21640 -14680
rect 22360 -14840 22380 -14680
rect 21620 -14860 22380 -14840
rect 23220 -14680 23980 -14610
rect 23220 -14840 23240 -14680
rect 23960 -14840 23980 -14680
rect 23220 -14860 23980 -14840
rect 25600 -14680 26400 -14660
rect 25600 -14840 25620 -14680
rect 26380 -14840 26400 -14680
rect 25600 -14910 26400 -14840
rect 27200 -14680 28000 -14660
rect 27200 -14840 27220 -14680
rect 27980 -14840 28000 -14680
rect 27200 -14910 28000 -14840
rect 32820 -14680 33580 -14610
rect 32820 -14840 32840 -14680
rect 33560 -14840 33580 -14680
rect 32820 -14860 33580 -14840
rect 36820 -14680 37580 -14610
rect 36820 -14840 36840 -14680
rect 37560 -14840 37580 -14680
rect 36820 -14860 37580 -14840
rect 39200 -14680 40000 -14660
rect 39200 -14840 39220 -14680
rect 39980 -14840 40000 -14680
rect 39200 -14910 40000 -14840
rect 40800 -14680 41600 -14660
rect 40800 -14840 40820 -14680
rect 41580 -14840 41600 -14680
rect 40800 -14910 41600 -14840
rect 42400 -14680 43200 -14660
rect 42400 -14840 42420 -14680
rect 43180 -14840 43200 -14680
rect 42400 -14910 43200 -14840
rect 44000 -14680 44800 -14660
rect 44000 -14840 44020 -14680
rect 44780 -14840 44800 -14680
rect 44000 -14910 44800 -14840
rect 46420 -14680 47180 -14610
rect 46420 -14840 46440 -14680
rect 47160 -14840 47180 -14680
rect 46420 -14860 47180 -14840
rect 14400 -15110 44800 -14910
<< viali >>
rect 41640 50 42360 3170
rect 41640 -4750 42360 -1630
rect -1560 -9790 -840 -6670
rect -760 -9790 -40 -6670
rect 8840 -9790 9560 -6670
rect 16840 -9790 17560 -6670
rect -1560 -14590 -840 -11470
rect -760 -14590 -40 -11470
rect 8840 -14590 9560 -11470
rect 13270 -9920 13310 -9880
rect 13270 -11380 13310 -11340
rect 21640 -9790 22360 -6670
rect 22440 -9790 23160 -6670
rect 41640 -9790 42360 -6670
rect 16840 -14590 17560 -11470
rect 21640 -14590 22360 -11470
rect 22440 -14590 23160 -11470
rect 41640 -14590 42360 -11470
<< metal1 >>
rect 41600 3170 42400 3210
rect 41600 50 41640 3170
rect 42360 50 42400 3170
rect 41600 -1630 42400 50
rect 41600 -4750 41640 -1630
rect 42360 -4750 42400 -1630
rect -1600 -6670 23200 -6650
rect -1600 -9790 -1560 -6670
rect -840 -9790 -760 -6670
rect -40 -9790 8840 -6670
rect 9560 -9790 16840 -6670
rect 17560 -9790 21640 -6670
rect 22360 -9790 22440 -6670
rect 23160 -9790 23200 -6670
rect -1600 -9880 23200 -9790
rect -1600 -9920 13270 -9880
rect 13310 -9920 23200 -9880
rect -1600 -11340 23200 -9920
rect -1600 -11380 13270 -11340
rect 13310 -11380 23200 -11340
rect -1600 -11470 23200 -11380
rect -1600 -14590 -1560 -11470
rect -840 -14590 -760 -11470
rect -40 -14590 8840 -11470
rect 9560 -14590 16840 -11470
rect 17560 -14590 21640 -11470
rect 22360 -14590 22440 -11470
rect 23160 -14590 23200 -11470
rect -1600 -14610 23200 -14590
rect 41600 -6670 42400 -4750
rect 41600 -9790 41640 -6670
rect 42360 -9790 42400 -6670
rect 41600 -11470 42400 -9790
rect 41600 -14590 41640 -11470
rect 42360 -14590 42400 -11470
rect 20000 -14620 20860 -14610
rect 41600 -14630 42400 -14590
<< end >>
