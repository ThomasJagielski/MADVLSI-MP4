magic
tech sky130A
timestamp 1617372252
<< nmos >>
rect 0 0 300 1600
rect 600 0 900 1600
rect 1200 0 1500 1600
rect 1800 0 2100 1600
rect 2400 0 2700 1600
rect 3000 0 3300 1600
rect 3600 0 3900 1600
rect 4200 0 4500 1600
rect 4800 0 5100 1600
rect 5400 0 5700 1600
rect 6000 0 6300 1600
rect 6600 0 6900 1600
rect 7200 0 7500 1600
rect 7800 0 8100 1600
rect 8400 0 8700 1600
rect 9000 0 9300 1600
rect 9600 0 9900 1600
rect 10200 0 10500 1600
rect 10800 0 11100 1600
rect 0 -2000 300 -400
rect 600 -2000 900 -400
rect 1200 -2000 1500 -400
rect 1800 -2000 2100 -400
rect 2400 -2000 2700 -400
rect 3000 -2000 3300 -400
rect 3600 -2000 3900 -400
rect 4200 -2000 4500 -400
rect 4800 -2000 5100 -400
rect 5400 -2000 5700 -400
rect 6000 -2000 6300 -400
rect 6600 -2000 6900 -400
rect 7200 -2000 7500 -400
rect 7800 -2000 8100 -400
rect 8400 -2000 8700 -400
rect 9000 -2000 9300 -400
rect 9600 -2000 9900 -400
rect 10200 -2000 10500 -400
rect 10800 -2000 11100 -400
rect 0 -4000 300 -2400
rect 600 -4000 900 -2400
rect 1200 -4000 1500 -2400
rect 1800 -4000 2100 -2400
rect 2400 -4000 2700 -2400
rect 3000 -4000 3300 -2400
rect 3600 -4000 3900 -2400
rect 4200 -4000 4500 -2400
rect 4800 -4000 5100 -2400
rect 5400 -4000 5700 -2400
rect 6000 -4000 6300 -2400
rect 6600 -4000 6900 -2400
rect 7200 -4000 7500 -2400
rect 7800 -4000 8100 -2400
rect 8400 -4000 8700 -2400
rect 9000 -4000 9300 -2400
rect 9600 -4000 9900 -2400
rect 10200 -4000 10500 -2400
rect 10800 -4000 11100 -2400
<< ndiff >>
rect -300 1585 0 1600
rect -300 15 -285 1585
rect -15 15 0 1585
rect -300 0 0 15
rect 300 1585 600 1600
rect 300 15 315 1585
rect 585 15 600 1585
rect 300 0 600 15
rect 900 1585 1200 1600
rect 900 15 915 1585
rect 1185 15 1200 1585
rect 900 0 1200 15
rect 1500 1585 1800 1600
rect 1500 15 1515 1585
rect 1785 15 1800 1585
rect 1500 0 1800 15
rect 2100 1585 2400 1600
rect 2100 15 2115 1585
rect 2385 15 2400 1585
rect 2100 0 2400 15
rect 2700 1585 3000 1600
rect 2700 15 2715 1585
rect 2985 15 3000 1585
rect 2700 0 3000 15
rect 3300 1585 3600 1600
rect 3300 15 3315 1585
rect 3585 15 3600 1585
rect 3300 0 3600 15
rect 3900 1585 4200 1600
rect 3900 15 3915 1585
rect 4185 15 4200 1585
rect 3900 0 4200 15
rect 4500 1585 4800 1600
rect 4500 15 4515 1585
rect 4785 15 4800 1585
rect 4500 0 4800 15
rect 5100 1585 5400 1600
rect 5100 15 5115 1585
rect 5385 15 5400 1585
rect 5100 0 5400 15
rect 5700 1585 6000 1600
rect 5700 15 5715 1585
rect 5985 15 6000 1585
rect 5700 0 6000 15
rect 6300 1585 6600 1600
rect 6300 15 6315 1585
rect 6585 15 6600 1585
rect 6300 0 6600 15
rect 6900 1585 7200 1600
rect 6900 15 6915 1585
rect 7185 15 7200 1585
rect 6900 0 7200 15
rect 7500 1585 7800 1600
rect 7500 15 7515 1585
rect 7785 15 7800 1585
rect 7500 0 7800 15
rect 8100 1585 8400 1600
rect 8100 15 8115 1585
rect 8385 15 8400 1585
rect 8100 0 8400 15
rect 8700 1585 9000 1600
rect 8700 15 8715 1585
rect 8985 15 9000 1585
rect 8700 0 9000 15
rect 9300 1585 9600 1600
rect 9300 15 9315 1585
rect 9585 15 9600 1585
rect 9300 0 9600 15
rect 9900 1585 10200 1600
rect 9900 15 9915 1585
rect 10185 15 10200 1585
rect 9900 0 10200 15
rect 10500 1585 10800 1600
rect 10500 15 10515 1585
rect 10785 15 10800 1585
rect 10500 0 10800 15
rect 11100 1585 11400 1600
rect 11100 15 11115 1585
rect 11385 15 11400 1585
rect 11100 0 11400 15
rect -300 -415 0 -400
rect -300 -1985 -285 -415
rect -15 -1985 0 -415
rect -300 -2000 0 -1985
rect 300 -415 600 -400
rect 300 -1985 315 -415
rect 585 -1985 600 -415
rect 300 -2000 600 -1985
rect 900 -415 1200 -400
rect 900 -1985 915 -415
rect 1185 -1985 1200 -415
rect 900 -2000 1200 -1985
rect 1500 -415 1800 -400
rect 1500 -1985 1515 -415
rect 1785 -1985 1800 -415
rect 1500 -2000 1800 -1985
rect 2100 -415 2400 -400
rect 2100 -1985 2115 -415
rect 2385 -1985 2400 -415
rect 2100 -2000 2400 -1985
rect 2700 -415 3000 -400
rect 2700 -1985 2715 -415
rect 2985 -1985 3000 -415
rect 2700 -2000 3000 -1985
rect 3300 -415 3600 -400
rect 3300 -1985 3315 -415
rect 3585 -1985 3600 -415
rect 3300 -2000 3600 -1985
rect 3900 -415 4200 -400
rect 3900 -1985 3915 -415
rect 4185 -1985 4200 -415
rect 3900 -2000 4200 -1985
rect 4500 -415 4800 -400
rect 4500 -1985 4515 -415
rect 4785 -1985 4800 -415
rect 4500 -2000 4800 -1985
rect 5100 -415 5400 -400
rect 5100 -1985 5115 -415
rect 5385 -1985 5400 -415
rect 5100 -2000 5400 -1985
rect 5700 -415 6000 -400
rect 5700 -1985 5715 -415
rect 5985 -1985 6000 -415
rect 5700 -2000 6000 -1985
rect 6300 -415 6600 -400
rect 6300 -1985 6315 -415
rect 6585 -1985 6600 -415
rect 6300 -2000 6600 -1985
rect 6900 -415 7200 -400
rect 6900 -1985 6915 -415
rect 7185 -1985 7200 -415
rect 6900 -2000 7200 -1985
rect 7500 -415 7800 -400
rect 7500 -1985 7515 -415
rect 7785 -1985 7800 -415
rect 7500 -2000 7800 -1985
rect 8100 -415 8400 -400
rect 8100 -1985 8115 -415
rect 8385 -1985 8400 -415
rect 8100 -2000 8400 -1985
rect 8700 -415 9000 -400
rect 8700 -1985 8715 -415
rect 8985 -1985 9000 -415
rect 8700 -2000 9000 -1985
rect 9300 -415 9600 -400
rect 9300 -1985 9315 -415
rect 9585 -1985 9600 -415
rect 9300 -2000 9600 -1985
rect 9900 -415 10200 -400
rect 9900 -1985 9915 -415
rect 10185 -1985 10200 -415
rect 9900 -2000 10200 -1985
rect 10500 -415 10800 -400
rect 10500 -1985 10515 -415
rect 10785 -1985 10800 -415
rect 10500 -2000 10800 -1985
rect 11100 -415 11400 -400
rect 11100 -1985 11115 -415
rect 11385 -1985 11400 -415
rect 11100 -2000 11400 -1985
rect -300 -2415 0 -2400
rect -300 -3985 -285 -2415
rect -15 -3985 0 -2415
rect -300 -4000 0 -3985
rect 300 -2415 600 -2400
rect 300 -3985 315 -2415
rect 585 -3985 600 -2415
rect 300 -4000 600 -3985
rect 900 -2415 1200 -2400
rect 900 -3985 915 -2415
rect 1185 -3985 1200 -2415
rect 900 -4000 1200 -3985
rect 1500 -2415 1800 -2400
rect 1500 -3985 1515 -2415
rect 1785 -3985 1800 -2415
rect 1500 -4000 1800 -3985
rect 2100 -2415 2400 -2400
rect 2100 -3985 2115 -2415
rect 2385 -3985 2400 -2415
rect 2100 -4000 2400 -3985
rect 2700 -2415 3000 -2400
rect 2700 -3985 2715 -2415
rect 2985 -3985 3000 -2415
rect 2700 -4000 3000 -3985
rect 3300 -2415 3600 -2400
rect 3300 -3985 3315 -2415
rect 3585 -3985 3600 -2415
rect 3300 -4000 3600 -3985
rect 3900 -2415 4200 -2400
rect 3900 -3985 3915 -2415
rect 4185 -3985 4200 -2415
rect 3900 -4000 4200 -3985
rect 4500 -2415 4800 -2400
rect 4500 -3985 4515 -2415
rect 4785 -3985 4800 -2415
rect 4500 -4000 4800 -3985
rect 5100 -2415 5400 -2400
rect 5100 -3985 5115 -2415
rect 5385 -3985 5400 -2415
rect 5100 -4000 5400 -3985
rect 5700 -2415 6000 -2400
rect 5700 -3985 5715 -2415
rect 5985 -3985 6000 -2415
rect 5700 -4000 6000 -3985
rect 6300 -2415 6600 -2400
rect 6300 -3985 6315 -2415
rect 6585 -3985 6600 -2415
rect 6300 -4000 6600 -3985
rect 6900 -2415 7200 -2400
rect 6900 -3985 6915 -2415
rect 7185 -3985 7200 -2415
rect 6900 -4000 7200 -3985
rect 7500 -2415 7800 -2400
rect 7500 -3985 7515 -2415
rect 7785 -3985 7800 -2415
rect 7500 -4000 7800 -3985
rect 8100 -2415 8400 -2400
rect 8100 -3985 8115 -2415
rect 8385 -3985 8400 -2415
rect 8100 -4000 8400 -3985
rect 8700 -2415 9000 -2400
rect 8700 -3985 8715 -2415
rect 8985 -3985 9000 -2415
rect 8700 -4000 9000 -3985
rect 9300 -2415 9600 -2400
rect 9300 -3985 9315 -2415
rect 9585 -3985 9600 -2415
rect 9300 -4000 9600 -3985
rect 9900 -2415 10200 -2400
rect 9900 -3985 9915 -2415
rect 10185 -3985 10200 -2415
rect 9900 -4000 10200 -3985
rect 10500 -2415 10800 -2400
rect 10500 -3985 10515 -2415
rect 10785 -3985 10800 -2415
rect 10500 -4000 10800 -3985
rect 11100 -2415 11400 -2400
rect 11100 -3985 11115 -2415
rect 11385 -3985 11400 -2415
rect 11100 -4000 11400 -3985
<< ndiffc >>
rect -285 15 -15 1585
rect 315 15 585 1585
rect 915 15 1185 1585
rect 1515 15 1785 1585
rect 2115 15 2385 1585
rect 2715 15 2985 1585
rect 3315 15 3585 1585
rect 3915 15 4185 1585
rect 4515 15 4785 1585
rect 5115 15 5385 1585
rect 5715 15 5985 1585
rect 6315 15 6585 1585
rect 6915 15 7185 1585
rect 7515 15 7785 1585
rect 8115 15 8385 1585
rect 8715 15 8985 1585
rect 9315 15 9585 1585
rect 9915 15 10185 1585
rect 10515 15 10785 1585
rect 11115 15 11385 1585
rect -285 -1985 -15 -415
rect 315 -1985 585 -415
rect 915 -1985 1185 -415
rect 1515 -1985 1785 -415
rect 2115 -1985 2385 -415
rect 2715 -1985 2985 -415
rect 3315 -1985 3585 -415
rect 3915 -1985 4185 -415
rect 4515 -1985 4785 -415
rect 5115 -1985 5385 -415
rect 5715 -1985 5985 -415
rect 6315 -1985 6585 -415
rect 6915 -1985 7185 -415
rect 7515 -1985 7785 -415
rect 8115 -1985 8385 -415
rect 8715 -1985 8985 -415
rect 9315 -1985 9585 -415
rect 9915 -1985 10185 -415
rect 10515 -1985 10785 -415
rect 11115 -1985 11385 -415
rect -285 -3985 -15 -2415
rect 315 -3985 585 -2415
rect 915 -3985 1185 -2415
rect 1515 -3985 1785 -2415
rect 2115 -3985 2385 -2415
rect 2715 -3985 2985 -2415
rect 3315 -3985 3585 -2415
rect 3915 -3985 4185 -2415
rect 4515 -3985 4785 -2415
rect 5115 -3985 5385 -2415
rect 5715 -3985 5985 -2415
rect 6315 -3985 6585 -2415
rect 6915 -3985 7185 -2415
rect 7515 -3985 7785 -2415
rect 8115 -3985 8385 -2415
rect 8715 -3985 8985 -2415
rect 9315 -3985 9585 -2415
rect 9915 -3985 10185 -2415
rect 10515 -3985 10785 -2415
rect 11115 -3985 11385 -2415
<< psubdiff >>
rect 2225 1665 2275 1680
rect 2225 1645 2240 1665
rect 2260 1645 2275 1665
rect 2825 1665 2875 1680
rect 2225 1630 2275 1645
rect 2825 1645 2840 1665
rect 2860 1645 2875 1665
rect 4625 1665 4675 1680
rect 2825 1630 2875 1645
rect 4625 1645 4640 1665
rect 4660 1645 4675 1665
rect 5225 1665 5275 1680
rect 4625 1630 4675 1645
rect 5225 1645 5240 1665
rect 5260 1645 5275 1665
rect 6425 1665 6475 1680
rect 5225 1630 5275 1645
rect 6425 1645 6440 1665
rect 6460 1645 6475 1665
rect 7625 1665 7675 1680
rect 6425 1630 6475 1645
rect 7625 1645 7640 1665
rect 7660 1645 7675 1665
rect 8825 1665 8875 1680
rect 7625 1630 7675 1645
rect 8825 1645 8840 1665
rect 8860 1645 8875 1665
rect 8825 1630 8875 1645
rect -600 1585 -300 1600
rect -600 15 -585 1585
rect -315 15 -300 1585
rect -600 0 -300 15
rect 11400 1585 11700 1600
rect 11400 15 11415 1585
rect 11685 15 11700 1585
rect 11400 0 11700 15
rect 2225 -235 2275 -220
rect 2225 -255 2240 -235
rect 2260 -255 2275 -235
rect 2225 -270 2275 -255
rect 4025 -235 4075 -220
rect 4025 -255 4040 -235
rect 4060 -255 4075 -235
rect 4025 -270 4075 -255
rect 5825 -235 5875 -220
rect 5825 -255 5840 -235
rect 5860 -255 5875 -235
rect 5825 -270 5875 -255
rect 8225 -235 8275 -220
rect 8225 -255 8240 -235
rect 8260 -255 8275 -235
rect 8225 -270 8275 -255
rect 9425 -235 9475 -220
rect 9425 -255 9440 -235
rect 9460 -255 9475 -235
rect 9425 -270 9475 -255
rect -600 -415 -300 -400
rect -600 -1985 -585 -415
rect -315 -1985 -300 -415
rect -600 -2000 -300 -1985
rect 11400 -415 11700 -400
rect 11400 -1985 11415 -415
rect 11685 -1985 11700 -415
rect 11400 -2000 11700 -1985
rect 1625 -2335 1675 -2320
rect 1625 -2355 1640 -2335
rect 1660 -2355 1675 -2335
rect 1625 -2370 1675 -2355
rect 4025 -2335 4075 -2320
rect 4025 -2355 4040 -2335
rect 4060 -2355 4075 -2335
rect 4025 -2370 4075 -2355
rect 5825 -2330 5875 -2315
rect 5825 -2350 5840 -2330
rect 5860 -2350 5875 -2330
rect 7625 -2330 7675 -2315
rect 5825 -2365 5875 -2350
rect 7625 -2350 7640 -2330
rect 7660 -2350 7675 -2330
rect 7625 -2365 7675 -2350
rect 9425 -2330 9475 -2315
rect 9425 -2350 9440 -2330
rect 9460 -2350 9475 -2330
rect 9425 -2365 9475 -2350
rect -600 -2415 -300 -2400
rect -600 -3985 -585 -2415
rect -315 -3985 -300 -2415
rect -600 -4000 -300 -3985
rect 11400 -2415 11700 -2400
rect 11400 -3985 11415 -2415
rect 11685 -3985 11700 -2415
rect 11400 -4000 11700 -3985
rect 2225 -4045 2275 -4030
rect 2225 -4065 2240 -4045
rect 2260 -4065 2275 -4045
rect 4025 -4045 4075 -4030
rect 2225 -4080 2275 -4065
rect 4025 -4065 4040 -4045
rect 4060 -4065 4075 -4045
rect 5825 -4045 5875 -4030
rect 4025 -4080 4075 -4065
rect 5825 -4065 5840 -4045
rect 5860 -4065 5875 -4045
rect 7625 -4045 7675 -4030
rect 5825 -4080 5875 -4065
rect 7625 -4065 7640 -4045
rect 7660 -4065 7675 -4045
rect 7625 -4080 7675 -4065
rect 9300 -4060 9350 -4045
rect 9300 -4080 9315 -4060
rect 9335 -4080 9350 -4060
rect 9300 -4095 9350 -4080
<< psubdiffcont >>
rect 2240 1645 2260 1665
rect 2840 1645 2860 1665
rect 4640 1645 4660 1665
rect 5240 1645 5260 1665
rect 6440 1645 6460 1665
rect 7640 1645 7660 1665
rect 8840 1645 8860 1665
rect -585 15 -315 1585
rect 11415 15 11685 1585
rect 2240 -255 2260 -235
rect 4040 -255 4060 -235
rect 5840 -255 5860 -235
rect 8240 -255 8260 -235
rect 9440 -255 9460 -235
rect -585 -1985 -315 -415
rect 11415 -1985 11685 -415
rect 1640 -2355 1660 -2335
rect 4040 -2355 4060 -2335
rect 5840 -2350 5860 -2330
rect 7640 -2350 7660 -2330
rect 9440 -2350 9460 -2330
rect -585 -3985 -315 -2415
rect 11415 -3985 11685 -2415
rect 2240 -4065 2260 -4045
rect 4040 -4065 4060 -4045
rect 5840 -4065 5860 -4045
rect 7640 -4065 7660 -4045
rect 9315 -4080 9335 -4060
<< poly >>
rect 9860 1685 9900 1695
rect -170 1645 -130 1655
rect -170 1630 -160 1645
rect -295 1625 -160 1630
rect -140 1630 -130 1645
rect 430 1645 470 1655
rect 430 1630 440 1645
rect -140 1625 440 1630
rect 460 1630 470 1645
rect 1200 1640 2225 1655
rect 460 1625 900 1630
rect -295 1615 900 1625
rect 0 1600 300 1615
rect 600 1600 900 1615
rect 1200 1600 1500 1640
rect 1800 1600 2100 1640
rect 2275 1640 2825 1655
rect 2875 1640 4625 1655
rect 2400 1600 2700 1615
rect 3000 1600 3300 1640
rect 3600 1600 3900 1615
rect 4200 1600 4500 1640
rect 4675 1640 5225 1655
rect 5275 1640 6425 1655
rect 4800 1600 5100 1615
rect 5400 1600 5700 1640
rect 6475 1640 7625 1655
rect 6000 1600 6300 1615
rect 6600 1600 6900 1640
rect 7675 1640 8825 1655
rect 9860 1665 9870 1685
rect 9890 1665 9900 1685
rect 9860 1655 9900 1665
rect 7200 1600 7500 1615
rect 7800 1600 8100 1640
rect 8875 1640 9900 1655
rect 8400 1600 8700 1615
rect 9000 1600 9300 1640
rect 9600 1600 9900 1640
rect 10620 1645 10660 1655
rect 10620 1630 10630 1645
rect 10200 1625 10630 1630
rect 10650 1630 10660 1645
rect 11230 1645 11270 1655
rect 11230 1630 11240 1645
rect 10650 1625 11240 1630
rect 11260 1630 11270 1645
rect 11260 1625 11395 1630
rect 10200 1615 11395 1625
rect 10200 1600 10500 1615
rect 10800 1600 11100 1615
rect 0 -15 300 0
rect 600 -15 900 0
rect 1200 -15 1500 0
rect 1800 -15 2100 0
rect 2400 -15 2700 0
rect 3000 -15 3300 0
rect 3600 -15 3900 0
rect 4200 -15 4500 0
rect 4800 -15 5100 0
rect 5400 -15 5700 0
rect 6000 -15 6300 0
rect 6600 -15 6900 0
rect 7200 -15 7500 0
rect 7800 -15 8100 0
rect 8400 -15 8700 0
rect 9000 -15 9300 0
rect 9600 -15 9900 0
rect 10200 -15 10500 0
rect 10800 -15 11100 0
rect 2530 -25 2570 -15
rect 2530 -45 2540 -25
rect 2560 -45 2570 -25
rect 2530 -55 2570 -45
rect 3730 -25 3770 -15
rect 3730 -45 3740 -25
rect 3760 -45 3770 -25
rect 3730 -55 3770 -45
rect 4930 -25 4970 -15
rect 4930 -45 4940 -25
rect 4960 -45 4970 -25
rect 4930 -55 4970 -45
rect 6130 -25 6170 -15
rect 6130 -45 6140 -25
rect 6160 -45 6170 -25
rect 6130 -55 6170 -45
rect 7330 -25 7370 -15
rect 7330 -45 7340 -25
rect 7360 -45 7370 -25
rect 7330 -55 7370 -45
rect 8530 -25 8570 -15
rect 8530 -45 8540 -25
rect 8560 -45 8570 -25
rect 8530 -55 8570 -45
rect 3600 -280 3900 -265
rect 3600 -330 3615 -280
rect 1200 -345 3615 -330
rect 3885 -330 3900 -280
rect 6600 -280 6900 -265
rect 6600 -330 6615 -280
rect 3885 -345 6615 -330
rect 6885 -330 6900 -280
rect 9150 -330 9165 -15
rect 6885 -345 9300 -330
rect -170 -355 -130 -345
rect -170 -370 -160 -355
rect -295 -375 -160 -370
rect -140 -370 -130 -355
rect 430 -355 470 -345
rect 430 -370 440 -355
rect -140 -375 440 -370
rect 460 -370 470 -355
rect 460 -375 900 -370
rect -295 -385 900 -375
rect 0 -400 300 -385
rect 600 -400 900 -385
rect 1200 -400 1500 -345
rect 1800 -400 2100 -345
rect 2400 -400 2700 -345
rect 3000 -400 3300 -345
rect 3730 -355 3770 -345
rect 3730 -375 3740 -355
rect 3760 -375 3770 -355
rect 3730 -385 3770 -375
rect 3600 -400 3900 -385
rect 4200 -400 4500 -345
rect 4800 -400 5100 -345
rect 5400 -400 5700 -345
rect 6000 -400 6300 -345
rect 6730 -355 6770 -345
rect 6730 -375 6740 -355
rect 6760 -375 6770 -355
rect 6730 -385 6770 -375
rect 6600 -400 6900 -385
rect 7200 -400 7500 -345
rect 7800 -400 8100 -345
rect 8400 -400 8700 -345
rect 9000 -400 9300 -345
rect 10030 -355 10070 -345
rect 10030 -370 10040 -355
rect 9600 -375 10040 -370
rect 10060 -370 10070 -355
rect 10630 -355 10670 -345
rect 10630 -370 10640 -355
rect 10060 -375 10640 -370
rect 10660 -370 10670 -355
rect 11230 -355 11270 -345
rect 11230 -370 11240 -355
rect 10660 -375 11240 -370
rect 11260 -370 11270 -355
rect 11260 -375 11395 -370
rect 9600 -385 11395 -375
rect 9600 -400 9900 -385
rect 10200 -400 10500 -385
rect 10800 -400 11100 -385
rect 0 -2015 300 -2000
rect 600 -2015 900 -2000
rect 1200 -2015 1500 -2000
rect 1800 -2015 2100 -2000
rect 2400 -2015 2700 -2000
rect 3000 -2015 3300 -2000
rect 3600 -2015 3900 -2000
rect 4200 -2015 4500 -2000
rect 4800 -2015 5100 -2000
rect 5400 -2015 5700 -2000
rect 6000 -2015 6300 -2000
rect 6600 -2015 6900 -2000
rect 7200 -2015 7500 -2000
rect 7800 -2015 8100 -2000
rect 8400 -2015 8700 -2000
rect 9000 -2015 9300 -2000
rect 9600 -2015 9900 -2000
rect 10200 -2015 10500 -2000
rect 10800 -2015 11100 -2000
rect 1735 -2025 1775 -2015
rect 1735 -2045 1745 -2025
rect 1765 -2045 1775 -2025
rect 1735 -2055 1775 -2045
rect 4630 -2025 4670 -2015
rect 4630 -2045 4640 -2025
rect 4660 -2045 4670 -2025
rect 4630 -2055 4670 -2045
rect 7525 -2025 7565 -2015
rect 7525 -2045 7535 -2025
rect 7555 -2045 7565 -2025
rect 7525 -2055 7565 -2045
rect 8725 -2025 8765 -2015
rect 8725 -2045 8735 -2025
rect 8755 -2045 8765 -2025
rect 8725 -2055 8765 -2045
rect 1735 -2335 1750 -2055
rect 1735 -2345 1775 -2335
rect 1735 -2365 1745 -2345
rect 1765 -2365 1775 -2345
rect 1735 -2375 1775 -2365
rect 4630 -2345 4645 -2055
rect 7525 -2295 7540 -2055
rect 7525 -2305 7565 -2295
rect 4630 -2355 4670 -2345
rect 4630 -2375 4640 -2355
rect 4660 -2375 4670 -2355
rect 7525 -2325 7535 -2305
rect 7555 -2325 7565 -2305
rect 7525 -2335 7565 -2325
rect 8725 -2340 8740 -2055
rect 8725 -2350 8765 -2340
rect 4630 -2385 4670 -2375
rect 8725 -2370 8735 -2350
rect 8755 -2370 8765 -2350
rect 8725 -2380 8765 -2370
rect 0 -2400 300 -2385
rect 600 -2400 900 -2385
rect 1200 -2400 1500 -2385
rect 1800 -2400 2100 -2385
rect 2400 -2400 2700 -2385
rect 3000 -2400 3300 -2385
rect 3600 -2400 3900 -2385
rect 4200 -2400 4500 -2385
rect 4800 -2400 5100 -2385
rect 5400 -2400 5700 -2385
rect 6000 -2400 6300 -2385
rect 6600 -2400 6900 -2385
rect 7200 -2400 7500 -2385
rect 7800 -2400 8100 -2385
rect 8400 -2400 8700 -2385
rect 9000 -2400 9300 -2385
rect 9600 -2400 9900 -2385
rect 10200 -2400 10500 -2385
rect 10800 -2400 11100 -2385
rect 0 -4015 300 -4000
rect 600 -4015 900 -4000
rect 1200 -4015 1500 -4000
rect 1800 -4015 2100 -4000
rect 2400 -4015 2700 -4000
rect 3000 -4015 3300 -4000
rect 3600 -4015 3900 -4000
rect 4200 -4015 4500 -4000
rect 4800 -4015 5100 -4000
rect 5400 -4015 5700 -4000
rect 6000 -4015 6300 -4000
rect 6600 -4015 6900 -4000
rect 7200 -4015 7500 -4000
rect 7800 -4015 8100 -4000
rect 8400 -4015 8700 -4000
rect 9000 -4015 9300 -4000
rect 9600 -4015 9900 -4000
rect 10200 -4015 10500 -4000
rect 10800 -4015 11100 -4000
rect -295 -4025 2100 -4015
rect -295 -4030 -160 -4025
rect -170 -4045 -160 -4030
rect -140 -4030 440 -4025
rect -140 -4045 -130 -4030
rect -170 -4055 -130 -4045
rect 430 -4045 440 -4030
rect 460 -4030 1040 -4025
rect 460 -4045 470 -4030
rect 430 -4055 470 -4045
rect 1030 -4045 1040 -4030
rect 1060 -4030 1640 -4025
rect 1060 -4045 1070 -4030
rect 1030 -4055 1070 -4045
rect 1630 -4045 1640 -4030
rect 1660 -4030 2100 -4025
rect 3130 -4025 3170 -4015
rect 1660 -4045 1670 -4030
rect 1630 -4055 1670 -4045
rect 3130 -4045 3140 -4025
rect 3160 -4045 3170 -4025
rect 3130 -4055 3170 -4045
rect 3730 -4025 3770 -4015
rect 3730 -4045 3740 -4025
rect 3760 -4045 3770 -4025
rect 4330 -4025 4370 -4015
rect 3730 -4055 3770 -4045
rect 4330 -4045 4340 -4025
rect 4360 -4045 4370 -4025
rect 4330 -4055 4370 -4045
rect 4930 -4025 4970 -4015
rect 4930 -4045 4940 -4025
rect 4960 -4045 4970 -4025
rect 4930 -4055 4970 -4045
rect 5530 -4025 5570 -4015
rect 5530 -4045 5540 -4025
rect 5560 -4045 5570 -4025
rect 6130 -4025 6170 -4015
rect 5530 -4055 5570 -4045
rect 6130 -4045 6140 -4025
rect 6160 -4045 6170 -4025
rect 6130 -4055 6170 -4045
rect 6730 -4025 6770 -4015
rect 6730 -4045 6740 -4025
rect 6760 -4045 6770 -4025
rect 6730 -4055 6770 -4045
rect 7330 -4025 7370 -4015
rect 7330 -4045 7340 -4025
rect 7360 -4045 7370 -4025
rect 7930 -4025 7970 -4015
rect 7330 -4055 7370 -4045
rect 7930 -4045 7940 -4025
rect 7960 -4045 7970 -4025
rect 8400 -4025 11395 -4015
rect 8400 -4030 8840 -4025
rect 7930 -4055 7970 -4045
rect 8830 -4045 8840 -4030
rect 8860 -4030 9440 -4025
rect 8860 -4045 8870 -4030
rect 9430 -4045 9440 -4030
rect 9460 -4030 10040 -4025
rect 9460 -4045 9470 -4030
rect 8830 -4055 8870 -4045
rect 9430 -4055 9470 -4045
rect 10030 -4045 10040 -4030
rect 10060 -4030 10640 -4025
rect 10060 -4045 10070 -4030
rect 10030 -4055 10070 -4045
rect 10630 -4045 10640 -4030
rect 10660 -4030 11240 -4025
rect 10660 -4045 10670 -4030
rect 10630 -4055 10670 -4045
rect 11230 -4045 11240 -4030
rect 11260 -4030 11395 -4025
rect 11260 -4045 11270 -4030
rect 11230 -4055 11270 -4045
<< polycont >>
rect -160 1625 -140 1645
rect 440 1625 460 1645
rect 9870 1665 9890 1685
rect 10630 1625 10650 1645
rect 11240 1625 11260 1645
rect 2540 -45 2560 -25
rect 3740 -45 3760 -25
rect 4940 -45 4960 -25
rect 6140 -45 6160 -25
rect 7340 -45 7360 -25
rect 8540 -45 8560 -25
rect -160 -375 -140 -355
rect 440 -375 460 -355
rect 3740 -375 3760 -355
rect 6740 -375 6760 -355
rect 10040 -375 10060 -355
rect 10640 -375 10660 -355
rect 11240 -375 11260 -355
rect 1745 -2045 1765 -2025
rect 4640 -2045 4660 -2025
rect 7535 -2045 7555 -2025
rect 8735 -2045 8755 -2025
rect 1745 -2365 1765 -2345
rect 4640 -2375 4660 -2355
rect 7535 -2325 7555 -2305
rect 8735 -2370 8755 -2350
rect -160 -4045 -140 -4025
rect 440 -4045 460 -4025
rect 1040 -4045 1060 -4025
rect 1640 -4045 1660 -4025
rect 3140 -4045 3160 -4025
rect 3740 -4045 3760 -4025
rect 4340 -4045 4360 -4025
rect 4940 -4045 4960 -4025
rect 5540 -4045 5560 -4025
rect 6140 -4045 6160 -4025
rect 6740 -4045 6760 -4025
rect 7340 -4045 7360 -4025
rect 7940 -4045 7960 -4025
rect 8840 -4045 8860 -4025
rect 9440 -4045 9460 -4025
rect 10040 -4045 10060 -4025
rect 10640 -4045 10660 -4025
rect 11240 -4045 11260 -4025
<< locali >>
rect 9305 1740 11700 1760
rect 2230 1710 2270 1720
rect 2230 1690 2240 1710
rect 2260 1690 2270 1710
rect 2230 1665 2270 1690
rect -170 1645 -130 1655
rect -170 1625 -160 1645
rect -140 1625 -130 1645
rect -170 1615 -130 1625
rect 430 1645 470 1655
rect 430 1625 440 1645
rect 460 1625 470 1645
rect 2230 1645 2240 1665
rect 2260 1645 2270 1665
rect 2230 1635 2270 1645
rect 2830 1710 2870 1720
rect 2830 1690 2840 1710
rect 2860 1690 2870 1710
rect 2830 1665 2870 1690
rect 2830 1645 2840 1665
rect 2860 1645 2870 1665
rect 2830 1635 2870 1645
rect 4630 1710 4670 1720
rect 4630 1690 4640 1710
rect 4660 1690 4670 1710
rect 4630 1665 4670 1690
rect 4630 1645 4640 1665
rect 4660 1645 4670 1665
rect 4630 1635 4670 1645
rect 5230 1710 5270 1720
rect 5230 1690 5240 1710
rect 5260 1690 5270 1710
rect 5230 1665 5270 1690
rect 5230 1645 5240 1665
rect 5260 1645 5270 1665
rect 5230 1635 5270 1645
rect 6430 1710 6470 1720
rect 6430 1690 6440 1710
rect 6460 1690 6470 1710
rect 6430 1665 6470 1690
rect 6430 1645 6440 1665
rect 6460 1645 6470 1665
rect 6430 1635 6470 1645
rect 7630 1710 7670 1720
rect 7630 1690 7640 1710
rect 7660 1690 7670 1710
rect 7630 1665 7670 1690
rect 7630 1645 7640 1665
rect 7660 1645 7670 1665
rect 7630 1635 7670 1645
rect 8830 1710 8870 1720
rect 8830 1690 8840 1710
rect 8860 1690 8870 1710
rect 8830 1665 8870 1690
rect 8830 1645 8840 1665
rect 8860 1645 8870 1665
rect 8830 1635 8870 1645
rect 430 1615 470 1625
rect -295 1595 -5 1615
rect -595 1585 -5 1595
rect -595 15 -585 1585
rect -315 15 -285 1585
rect -15 15 -5 1585
rect -595 5 -5 15
rect 305 1585 595 1615
rect 305 15 315 1585
rect 585 15 595 1585
rect 305 5 595 15
rect 905 1585 1195 1595
rect 905 15 915 1585
rect 1185 15 1195 1585
rect 905 -20 1195 15
rect 1505 1585 1795 1595
rect 1505 15 1515 1585
rect 1785 15 1795 1585
rect 1505 5 1795 15
rect 2105 1585 2400 1595
rect 2105 15 2115 1585
rect 2385 15 2400 1585
rect 2105 5 2400 15
rect 2705 1585 2995 1595
rect 2705 15 2715 1585
rect 2985 15 2995 1585
rect 2105 -20 2395 5
rect 905 -40 2395 -20
rect 2530 -25 2570 -15
rect -170 -355 -130 -345
rect -170 -375 -160 -355
rect -140 -375 -130 -355
rect -170 -385 -130 -375
rect 430 -355 470 -345
rect 430 -375 440 -355
rect 460 -375 470 -355
rect 430 -385 470 -375
rect 1640 -385 1660 -40
rect 2530 -45 2540 -25
rect 2560 -45 2570 -25
rect 2705 -40 2995 15
rect 3305 1585 3595 1595
rect 3305 15 3315 1585
rect 3585 15 3595 1585
rect 3305 5 3595 15
rect 3905 1585 4195 1595
rect 3905 15 3915 1585
rect 4185 15 4195 1585
rect 3905 5 4195 15
rect 4505 1585 4795 1595
rect 4505 15 4515 1585
rect 4785 15 4795 1585
rect 3730 -25 3770 -15
rect 2530 -65 2570 -45
rect 2530 -85 2540 -65
rect 2560 -85 2570 -65
rect 2530 -95 2570 -85
rect 2230 -190 2270 -180
rect 2230 -210 2240 -190
rect 2260 -210 2270 -190
rect 2230 -235 2270 -210
rect 2230 -255 2240 -235
rect 2260 -255 2270 -235
rect 2230 -265 2270 -255
rect 2840 -295 2860 -40
rect 3730 -45 3740 -25
rect 3760 -45 3770 -25
rect 4505 -40 4795 15
rect 5105 1585 5395 1595
rect 5105 15 5115 1585
rect 5385 15 5395 1585
rect 4930 -25 4970 -15
rect 3730 -65 3770 -45
rect 3730 -85 3740 -65
rect 3760 -85 3770 -65
rect 3730 -95 3770 -85
rect 4030 -190 4070 -180
rect 4030 -210 4040 -190
rect 4060 -210 4070 -190
rect 4030 -235 4070 -210
rect 4030 -255 4040 -235
rect 4060 -255 4070 -235
rect 2105 -315 2860 -295
rect 3600 -280 3900 -260
rect 4030 -265 4070 -255
rect -295 -405 -5 -385
rect -595 -415 -5 -405
rect -595 -1985 -585 -415
rect -315 -1985 -285 -415
rect -15 -1985 -5 -415
rect -595 -1995 -5 -1985
rect 305 -415 595 -385
rect 305 -1985 315 -415
rect 585 -1985 595 -415
rect 305 -1995 595 -1985
rect 905 -415 1195 -405
rect 905 -1985 915 -415
rect 1185 -1985 1195 -415
rect 905 -2080 1195 -1985
rect 1505 -415 1795 -385
rect 1505 -1985 1515 -415
rect 1785 -1985 1795 -415
rect 1505 -2015 1795 -1985
rect 2105 -405 2395 -315
rect 3600 -340 3620 -280
rect 2705 -360 3620 -340
rect 3730 -315 3770 -305
rect 3730 -335 3740 -315
rect 3760 -335 3770 -315
rect 3730 -355 3770 -335
rect 2105 -415 2400 -405
rect 2105 -1985 2115 -415
rect 2385 -1985 2400 -415
rect 2105 -1995 2400 -1985
rect 2705 -415 2995 -360
rect 3730 -375 3740 -355
rect 3760 -375 3770 -355
rect 3880 -340 3900 -280
rect 4640 -340 4660 -40
rect 4930 -45 4940 -25
rect 4960 -45 4970 -25
rect 5105 -35 5395 15
rect 5705 1585 5995 1595
rect 5705 15 5715 1585
rect 5985 15 5995 1585
rect 5705 5 5995 15
rect 6305 1585 6595 1595
rect 6305 15 6315 1585
rect 6585 15 6595 1585
rect 6130 -25 6170 -15
rect 4930 -65 4970 -45
rect 4930 -85 4940 -65
rect 4960 -85 4970 -65
rect 4930 -95 4970 -85
rect 5240 -340 5260 -35
rect 6130 -45 6140 -25
rect 6160 -45 6170 -25
rect 6305 -35 6595 15
rect 6905 1585 7195 1595
rect 6905 15 6915 1585
rect 7185 15 7195 1585
rect 6905 5 7195 15
rect 7505 1585 7795 1595
rect 7505 15 7515 1585
rect 7785 15 7795 1585
rect 6130 -65 6170 -45
rect 6130 -85 6140 -65
rect 6160 -85 6170 -65
rect 6130 -95 6170 -85
rect 5830 -190 5870 -180
rect 5830 -210 5840 -190
rect 5860 -210 5870 -190
rect 5830 -235 5870 -210
rect 5830 -255 5840 -235
rect 5860 -255 5870 -235
rect 5830 -265 5870 -255
rect 6575 -260 6595 -35
rect 7330 -25 7370 -15
rect 7330 -45 7340 -25
rect 7360 -45 7370 -25
rect 7505 -35 7795 15
rect 8105 1585 8395 1595
rect 8105 15 8115 1585
rect 8385 15 8395 1585
rect 8105 5 8395 15
rect 8705 1585 8995 1595
rect 8705 15 8715 1585
rect 8985 15 8995 1585
rect 8530 -25 8570 -15
rect 7330 -65 7370 -45
rect 7330 -85 7340 -65
rect 7360 -85 7370 -65
rect 7330 -95 7370 -85
rect 6575 -280 6900 -260
rect 6730 -315 6770 -305
rect 6730 -335 6740 -315
rect 6760 -335 6770 -315
rect 3880 -360 4795 -340
rect 3730 -385 3770 -375
rect 2705 -1985 2715 -415
rect 2985 -1985 2995 -415
rect 2705 -1995 2995 -1985
rect 3305 -415 3595 -405
rect 3305 -1985 3315 -415
rect 3585 -1985 3595 -415
rect 1735 -2025 1775 -2015
rect 1735 -2045 1745 -2025
rect 1765 -2045 1775 -2025
rect 1735 -2055 1775 -2045
rect 2105 -2080 2395 -1995
rect 3305 -2080 3595 -1985
rect 905 -2100 3595 -2080
rect 3905 -415 4195 -405
rect 3905 -1985 3915 -415
rect 4185 -1985 4195 -415
rect 3905 -2080 4195 -1985
rect 4505 -415 4795 -360
rect 4505 -1985 4515 -415
rect 4785 -1985 4795 -415
rect 4505 -2015 4795 -1985
rect 5105 -360 6325 -340
rect 5105 -415 5395 -360
rect 6305 -385 6325 -360
rect 6730 -355 6770 -335
rect 6730 -375 6740 -355
rect 6760 -375 6770 -355
rect 6880 -340 6900 -280
rect 7640 -295 7660 -35
rect 8530 -45 8540 -25
rect 8560 -45 8570 -25
rect 8705 -20 8995 15
rect 9305 1585 9595 1740
rect 9860 1685 11700 1695
rect 9860 1665 9870 1685
rect 9890 1675 11700 1685
rect 9890 1665 9900 1675
rect 9860 1655 9900 1665
rect 10620 1645 10660 1655
rect 10620 1625 10630 1645
rect 10650 1625 10660 1645
rect 10620 1615 10660 1625
rect 11230 1645 11270 1655
rect 11230 1625 11240 1645
rect 11260 1625 11270 1645
rect 11230 1615 11270 1625
rect 9305 15 9315 1585
rect 9585 15 9595 1585
rect 9305 5 9595 15
rect 9905 1585 10195 1595
rect 9905 15 9915 1585
rect 10185 15 10195 1585
rect 9905 -20 10195 15
rect 10505 1585 10795 1615
rect 10505 15 10515 1585
rect 10785 15 10795 1585
rect 10505 5 10795 15
rect 11105 1595 11395 1615
rect 11105 1585 11695 1595
rect 11105 15 11115 1585
rect 11385 15 11415 1585
rect 11685 15 11695 1585
rect 11105 5 11695 15
rect 8705 -40 10195 -20
rect 8530 -65 8570 -45
rect 8530 -85 8540 -65
rect 8560 -85 8570 -65
rect 8530 -95 8570 -85
rect 8230 -190 8270 -180
rect 8230 -210 8240 -190
rect 8260 -210 8270 -190
rect 8230 -235 8270 -210
rect 8230 -255 8240 -235
rect 8260 -255 8270 -235
rect 8230 -265 8270 -255
rect 7640 -315 8395 -295
rect 6880 -360 7795 -340
rect 6730 -385 6770 -375
rect 5105 -1985 5115 -415
rect 5385 -1985 5395 -415
rect 4630 -2025 4670 -2015
rect 4630 -2045 4640 -2025
rect 4660 -2045 4670 -2025
rect 4630 -2055 4670 -2045
rect 5105 -2080 5395 -1985
rect 5705 -415 5995 -405
rect 5705 -1985 5715 -415
rect 5985 -1985 5995 -415
rect 5705 -2015 5995 -1985
rect 6305 -415 6595 -385
rect 6305 -1985 6315 -415
rect 6585 -1985 6595 -415
rect 6305 -1995 6595 -1985
rect 6905 -415 7195 -405
rect 6905 -1985 6915 -415
rect 7185 -1985 7195 -415
rect 3905 -2100 5395 -2080
rect 1630 -2335 1670 -2325
rect 1630 -2355 1640 -2335
rect 1660 -2355 1670 -2335
rect 1630 -2405 1670 -2355
rect 1735 -2345 1775 -2335
rect 1735 -2365 1745 -2345
rect 1765 -2355 1775 -2345
rect 1765 -2365 2995 -2355
rect 1735 -2375 2995 -2365
rect -595 -2415 -5 -2405
rect -595 -3985 -585 -2415
rect -315 -3985 -285 -2415
rect -15 -3985 -5 -2415
rect -595 -3995 -5 -3985
rect -295 -4015 -5 -3995
rect 305 -2415 595 -2405
rect 305 -3985 315 -2415
rect 585 -3985 595 -2415
rect 305 -4015 595 -3985
rect 905 -2415 1195 -2405
rect 905 -3985 915 -2415
rect 1185 -3985 1195 -2415
rect 905 -4015 1195 -3985
rect 1505 -2415 1795 -2405
rect 1505 -3985 1515 -2415
rect 1785 -3985 1795 -2415
rect 1505 -4015 1795 -3985
rect 2105 -2415 2400 -2405
rect 2105 -3985 2115 -2415
rect 2385 -3985 2400 -2415
rect 2105 -3995 2400 -3985
rect 2705 -2415 2995 -2375
rect 3440 -2385 3460 -2100
rect 4030 -2335 4070 -2325
rect 4030 -2355 4040 -2335
rect 4060 -2355 4070 -2335
rect 2705 -3985 2715 -2415
rect 2985 -3985 2995 -2415
rect 2705 -3995 2995 -3985
rect 3305 -2415 3595 -2385
rect 4030 -2405 4070 -2355
rect 4630 -2355 4670 -2345
rect 4630 -2375 4640 -2355
rect 4660 -2375 4670 -2355
rect 4630 -2385 4670 -2375
rect 5240 -2385 5260 -2100
rect 5975 -2315 5995 -2015
rect 6905 -2080 7195 -1985
rect 7505 -415 7795 -360
rect 7505 -1985 7515 -415
rect 7785 -1985 7795 -415
rect 7505 -2015 7795 -1985
rect 8105 -415 8395 -315
rect 8840 -390 8860 -40
rect 9430 -190 9470 -180
rect 9430 -210 9440 -190
rect 9460 -210 9470 -190
rect 9430 -235 9470 -210
rect 9430 -255 9440 -235
rect 9460 -255 9470 -235
rect 9430 -265 9470 -255
rect 10030 -355 10070 -345
rect 10030 -375 10040 -355
rect 10060 -375 10070 -355
rect 10030 -385 10070 -375
rect 10630 -355 10670 -345
rect 10630 -375 10640 -355
rect 10660 -375 10670 -355
rect 10630 -385 10670 -375
rect 11230 -355 11270 -345
rect 11230 -375 11240 -355
rect 11260 -375 11270 -355
rect 11230 -385 11270 -375
rect 8105 -1985 8115 -415
rect 8385 -1985 8395 -415
rect 7525 -2025 7565 -2015
rect 7525 -2045 7535 -2025
rect 7555 -2045 7565 -2025
rect 7525 -2055 7565 -2045
rect 8105 -2080 8395 -1985
rect 8705 -415 8995 -390
rect 8705 -1985 8715 -415
rect 8985 -1985 8995 -415
rect 8705 -2015 8995 -1985
rect 9305 -415 9595 -405
rect 9305 -1985 9315 -415
rect 9585 -1985 9595 -415
rect 8725 -2025 8765 -2015
rect 8725 -2045 8735 -2025
rect 8755 -2045 8765 -2025
rect 8725 -2055 8765 -2045
rect 9305 -2080 9595 -1985
rect 9905 -415 10195 -385
rect 9905 -1985 9915 -415
rect 10185 -1985 10195 -415
rect 9905 -1995 10195 -1985
rect 10505 -415 10795 -385
rect 10505 -1985 10515 -415
rect 10785 -1985 10795 -415
rect 10505 -1995 10795 -1985
rect 11105 -405 11395 -385
rect 11105 -415 11695 -405
rect 11105 -1985 11115 -415
rect 11385 -1985 11415 -415
rect 11685 -1985 11695 -415
rect 11105 -1995 11695 -1985
rect 6905 -2100 9595 -2080
rect 7525 -2305 7565 -2295
rect 7525 -2315 7535 -2305
rect 5830 -2330 5870 -2320
rect 5830 -2350 5840 -2330
rect 5860 -2350 5870 -2330
rect 5975 -2325 7535 -2315
rect 7555 -2325 7565 -2305
rect 5975 -2335 7565 -2325
rect 3305 -3985 3315 -2415
rect 3585 -3985 3595 -2415
rect 3305 -3995 3595 -3985
rect 3905 -2415 4195 -2405
rect 3905 -3985 3915 -2415
rect 4185 -3985 4195 -2415
rect 3905 -3995 4195 -3985
rect 4505 -2415 4795 -2385
rect 4505 -3985 4515 -2415
rect 4785 -3985 4795 -2415
rect 4505 -3995 4795 -3985
rect 5105 -2415 5395 -2385
rect 5830 -2405 5870 -2350
rect 5105 -3985 5115 -2415
rect 5385 -3985 5395 -2415
rect 5105 -3995 5395 -3985
rect 5705 -2415 5995 -2405
rect 5705 -3985 5715 -2415
rect 5985 -3985 5995 -2415
rect 5705 -3995 5995 -3985
rect 6305 -2415 6595 -2335
rect 7590 -2360 7610 -2100
rect 6305 -3985 6315 -2415
rect 6585 -3985 6595 -2415
rect 6305 -3995 6595 -3985
rect 6905 -2380 7610 -2360
rect 7630 -2330 7670 -2320
rect 7630 -2350 7640 -2330
rect 7660 -2350 7670 -2330
rect 9430 -2330 9470 -2320
rect 6905 -2415 7195 -2380
rect 7630 -2405 7670 -2350
rect 8725 -2350 8765 -2340
rect 8725 -2360 8735 -2350
rect 8105 -2370 8735 -2360
rect 8755 -2370 8765 -2350
rect 8105 -2380 8765 -2370
rect 9430 -2350 9440 -2330
rect 9460 -2350 9470 -2330
rect 6905 -3985 6915 -2415
rect 7185 -3985 7195 -2415
rect 6905 -3995 7195 -3985
rect 7505 -2415 7795 -2405
rect 7505 -3985 7515 -2415
rect 7785 -3985 7795 -2415
rect 7505 -3995 7795 -3985
rect 8105 -2415 8395 -2380
rect 9430 -2405 9470 -2350
rect 8105 -3985 8115 -2415
rect 8385 -3985 8395 -2415
rect 8105 -3995 8395 -3985
rect 8705 -2415 8995 -2405
rect 8705 -3985 8715 -2415
rect 8985 -3985 8995 -2415
rect -170 -4025 -130 -4015
rect -170 -4045 -160 -4025
rect -140 -4045 -130 -4025
rect -170 -4055 -130 -4045
rect 430 -4025 470 -4015
rect 430 -4045 440 -4025
rect 460 -4045 470 -4025
rect 430 -4055 470 -4045
rect 1030 -4025 1070 -4015
rect 1030 -4045 1040 -4025
rect 1060 -4045 1070 -4025
rect 1030 -4055 1070 -4045
rect 1630 -4025 1670 -4015
rect 1630 -4045 1640 -4025
rect 1660 -4045 1670 -4025
rect 1630 -4055 1670 -4045
rect 2230 -4045 2270 -3995
rect 2230 -4065 2240 -4045
rect 2260 -4065 2270 -4045
rect 2230 -4075 2270 -4065
rect 3130 -4025 3170 -4015
rect 3130 -4045 3140 -4025
rect 3160 -4045 3170 -4025
rect 3130 -4090 3170 -4045
rect 3130 -4110 3140 -4090
rect 3160 -4110 3170 -4090
rect 3730 -4025 3770 -4015
rect 3730 -4045 3740 -4025
rect 3760 -4045 3770 -4025
rect 3730 -4065 3770 -4045
rect 3730 -4085 3740 -4065
rect 3760 -4085 3770 -4065
rect 4030 -4045 4070 -3995
rect 4030 -4065 4040 -4045
rect 4060 -4065 4070 -4045
rect 4030 -4075 4070 -4065
rect 4330 -4025 4370 -4015
rect 4330 -4045 4340 -4025
rect 4360 -4045 4370 -4025
rect 3730 -4095 3770 -4085
rect 4330 -4090 4370 -4045
rect 3130 -4120 3170 -4110
rect 4330 -4110 4340 -4090
rect 4360 -4110 4370 -4090
rect 4330 -4120 4370 -4110
rect 4930 -4025 4970 -4015
rect 4930 -4045 4940 -4025
rect 4960 -4045 4970 -4025
rect 4930 -4090 4970 -4045
rect 4930 -4110 4940 -4090
rect 4960 -4110 4970 -4090
rect 4930 -4120 4970 -4110
rect 5530 -4025 5570 -4015
rect 5530 -4045 5540 -4025
rect 5560 -4045 5570 -4025
rect 5530 -4090 5570 -4045
rect 5830 -4045 5870 -3995
rect 5830 -4065 5840 -4045
rect 5860 -4065 5870 -4045
rect 5830 -4075 5870 -4065
rect 6130 -4025 6170 -4015
rect 6130 -4045 6140 -4025
rect 6160 -4045 6170 -4025
rect 5530 -4110 5540 -4090
rect 5560 -4110 5570 -4090
rect 5530 -4120 5570 -4110
rect 6130 -4090 6170 -4045
rect 6130 -4110 6140 -4090
rect 6160 -4110 6170 -4090
rect 6130 -4120 6170 -4110
rect 6730 -4025 6770 -4015
rect 6730 -4045 6740 -4025
rect 6760 -4045 6770 -4025
rect 6730 -4090 6770 -4045
rect 6730 -4110 6740 -4090
rect 6760 -4110 6770 -4090
rect 6730 -4120 6770 -4110
rect 7330 -4025 7370 -4015
rect 7330 -4045 7340 -4025
rect 7360 -4045 7370 -4025
rect 7330 -4090 7370 -4045
rect 7630 -4045 7670 -3995
rect 8705 -4015 8995 -3985
rect 9305 -2415 9595 -2405
rect 9305 -3985 9315 -2415
rect 9585 -3985 9595 -2415
rect 9305 -4015 9595 -3985
rect 9905 -2415 10195 -2405
rect 9905 -3985 9915 -2415
rect 10185 -3985 10195 -2415
rect 9905 -4015 10195 -3985
rect 10505 -2415 10795 -2405
rect 10505 -3985 10515 -2415
rect 10785 -3985 10795 -2415
rect 10505 -4015 10795 -3985
rect 11105 -2415 11695 -2405
rect 11105 -3985 11115 -2415
rect 11385 -3985 11415 -2415
rect 11685 -3985 11695 -2415
rect 11105 -3995 11695 -3985
rect 11105 -4015 11395 -3995
rect 7630 -4065 7640 -4045
rect 7660 -4065 7670 -4045
rect 7630 -4075 7670 -4065
rect 7930 -4025 7970 -4015
rect 7930 -4045 7940 -4025
rect 7960 -4045 7970 -4025
rect 7330 -4110 7340 -4090
rect 7360 -4110 7370 -4090
rect 7330 -4120 7370 -4110
rect 7930 -4090 7970 -4045
rect 8830 -4025 8870 -4015
rect 8830 -4045 8840 -4025
rect 8860 -4045 8870 -4025
rect 8830 -4055 8870 -4045
rect 9305 -4060 9345 -4015
rect 9430 -4025 9470 -4015
rect 9430 -4045 9440 -4025
rect 9460 -4045 9470 -4025
rect 9430 -4055 9470 -4045
rect 10030 -4025 10070 -4015
rect 10030 -4045 10040 -4025
rect 10060 -4045 10070 -4025
rect 10030 -4055 10070 -4045
rect 10630 -4025 10670 -4015
rect 10630 -4045 10640 -4025
rect 10660 -4045 10670 -4025
rect 10630 -4055 10670 -4045
rect 11230 -4025 11270 -4015
rect 11230 -4045 11240 -4025
rect 11260 -4045 11270 -4025
rect 11230 -4055 11270 -4045
rect 9305 -4080 9315 -4060
rect 9335 -4080 9345 -4060
rect 9305 -4090 9345 -4080
rect 7930 -4110 7940 -4090
rect 7960 -4110 7970 -4090
rect 7930 -4120 7970 -4110
<< viali >>
rect 2240 1690 2260 1710
rect 2840 1690 2860 1710
rect 4640 1690 4660 1710
rect 5240 1690 5260 1710
rect 6440 1690 6460 1710
rect 7640 1690 7660 1710
rect 8840 1690 8860 1710
rect -585 15 -315 1585
rect -285 15 -15 1585
rect 315 15 585 1585
rect 1515 15 1785 1585
rect 3315 15 3585 1585
rect 3915 15 4185 1585
rect 2540 -85 2560 -65
rect 2240 -210 2260 -190
rect 3740 -85 3760 -65
rect 4040 -210 4060 -190
rect -585 -1985 -315 -415
rect -285 -1985 -15 -415
rect 315 -1985 585 -415
rect 3740 -335 3760 -315
rect 5715 15 5985 1585
rect 4940 -85 4960 -65
rect 6915 15 7185 1585
rect 6140 -85 6160 -65
rect 5840 -210 5860 -190
rect 8115 15 8385 1585
rect 7340 -85 7360 -65
rect 6740 -335 6760 -315
rect 10515 15 10785 1585
rect 11115 15 11385 1585
rect 11415 15 11685 1585
rect 8540 -85 8560 -65
rect 8240 -210 8260 -190
rect -585 -3985 -315 -2415
rect -285 -3985 -15 -2415
rect 315 -3985 585 -2415
rect 915 -3985 1185 -2415
rect 1515 -3985 1785 -2415
rect 2115 -3985 2385 -2415
rect 9440 -210 9460 -190
rect 9915 -1985 10185 -415
rect 10515 -1985 10785 -415
rect 11115 -1985 11385 -415
rect 11415 -1985 11685 -415
rect 3915 -3985 4185 -2415
rect 5715 -3985 5985 -2415
rect 7515 -3985 7785 -2415
rect 8715 -3985 8985 -2415
rect 3140 -4110 3160 -4090
rect 3740 -4085 3760 -4065
rect 4340 -4110 4360 -4090
rect 4940 -4110 4960 -4090
rect 5540 -4110 5560 -4090
rect 6140 -4110 6160 -4090
rect 6740 -4110 6760 -4090
rect 9315 -3985 9585 -2415
rect 9915 -3985 10185 -2415
rect 10515 -3985 10785 -2415
rect 11115 -3985 11385 -2415
rect 11415 -3985 11685 -2415
rect 7340 -4110 7360 -4090
rect 7940 -4110 7960 -4090
<< metal1 >>
rect -600 1815 11700 3405
rect -600 1585 595 1595
rect -600 15 -585 1585
rect -315 15 -285 1585
rect -15 15 315 1585
rect 585 15 595 1585
rect -600 -400 595 15
rect 1505 1585 1795 1815
rect 1505 15 1515 1585
rect 1785 15 1795 1585
rect 1505 5 1795 15
rect 2105 1710 2395 1730
rect 2105 1690 2240 1710
rect 2260 1690 2395 1710
rect 2105 -190 2395 1690
rect 2705 1710 2995 1730
rect 2705 1690 2840 1710
rect 2860 1690 2995 1710
rect 2105 -210 2240 -190
rect 2260 -210 2395 -190
rect 2105 -400 2395 -210
rect 2530 -65 2570 -55
rect 2530 -85 2540 -65
rect 2560 -85 2570 -65
rect 2530 -400 2570 -85
rect 2705 -400 2995 1690
rect 3305 1585 3595 1815
rect 3305 15 3315 1585
rect 3585 15 3595 1585
rect 3305 5 3595 15
rect 3905 1585 4195 1815
rect 4505 1710 4795 1730
rect 4505 1690 4640 1710
rect 4660 1690 4795 1710
rect 4505 1600 4795 1690
rect 5105 1710 5395 1730
rect 5105 1690 5240 1710
rect 5260 1690 5395 1710
rect 5105 1600 5395 1690
rect 3905 15 3915 1585
rect 4185 15 4195 1585
rect 5705 1585 5995 1815
rect 3905 5 4195 15
rect 3730 -65 3770 -15
rect 3730 -85 3740 -65
rect 3760 -85 3770 -65
rect 3730 -315 3770 -85
rect 3730 -335 3740 -315
rect 3760 -335 3770 -315
rect 3730 -400 3770 -335
rect 3905 -190 4195 -170
rect 3905 -210 4040 -190
rect 4060 -210 4195 -190
rect 3905 -400 4195 -210
rect 4505 -400 4795 1565
rect 4930 -65 4970 -15
rect 4930 -85 4940 -65
rect 4960 -85 4970 -65
rect 4930 -400 4970 -85
rect 5105 -400 5395 1570
rect 5705 15 5715 1585
rect 5985 15 5995 1585
rect 5705 5 5995 15
rect 6305 1710 6595 1730
rect 6305 1690 6440 1710
rect 6460 1690 6595 1710
rect 6130 -65 6170 -15
rect 6130 -85 6140 -65
rect 6160 -85 6170 -65
rect 5705 -190 5995 -175
rect 5705 -210 5840 -190
rect 5860 -210 5995 -190
rect 5705 -400 5995 -210
rect 6130 -400 6170 -85
rect 6305 -400 6595 1690
rect 6905 1585 7195 1815
rect 6905 15 6915 1585
rect 7185 15 7195 1585
rect 6905 5 7195 15
rect 7505 1710 7795 1730
rect 7505 1690 7640 1710
rect 7660 1690 7795 1710
rect 7330 -65 7370 -15
rect 7330 -85 7340 -65
rect 7360 -85 7370 -65
rect 6730 -315 6770 -305
rect 6730 -335 6740 -315
rect 6760 -335 6770 -315
rect 6730 -400 6770 -335
rect 7330 -400 7370 -85
rect 7505 -400 7795 1690
rect 8105 1585 8395 1815
rect 8105 15 8115 1585
rect 8385 15 8395 1585
rect 8105 5 8395 15
rect 8705 1710 8995 1730
rect 8705 1690 8840 1710
rect 8860 1690 8995 1710
rect 8530 -65 8570 -15
rect 8530 -85 8540 -65
rect 8560 -85 8570 -65
rect 8105 -190 8395 -170
rect 8105 -210 8240 -190
rect 8260 -210 8395 -190
rect 8105 -400 8395 -210
rect 8530 -400 8570 -85
rect 8705 -400 8995 1690
rect 10505 1585 11695 1595
rect 10505 15 10515 1585
rect 10785 15 11115 1585
rect 11385 15 11415 1585
rect 11685 15 11695 1585
rect 9305 -190 9595 -175
rect 9305 -210 9440 -190
rect 9460 -210 9595 -190
rect 9305 -400 9595 -210
rect 10505 -400 11695 15
rect -600 -415 11700 -400
rect -600 -1985 -585 -415
rect -315 -1985 -285 -415
rect -15 -1985 315 -415
rect 585 -1985 9915 -415
rect 10185 -1985 10515 -415
rect 10785 -1985 11115 -415
rect 11385 -1985 11415 -415
rect 11685 -1985 11700 -415
rect -600 -2415 11700 -1985
rect -600 -3985 -585 -2415
rect -315 -3985 -285 -2415
rect -15 -3985 315 -2415
rect 585 -3985 915 -2415
rect 1185 -3985 1515 -2415
rect 1785 -3985 2115 -2415
rect 2385 -3985 3915 -2415
rect 4185 -3985 5715 -2415
rect 5985 -3985 7515 -2415
rect 7785 -3985 8715 -2415
rect 8985 -3985 9315 -2415
rect 9585 -3985 9915 -2415
rect 10185 -3985 10515 -2415
rect 10785 -3985 11115 -2415
rect 11385 -3985 11415 -2415
rect 11685 -3985 11700 -2415
rect -600 -3995 11700 -3985
rect 3130 -4090 3170 -3995
rect 3130 -4110 3140 -4090
rect 3160 -4110 3170 -4090
rect 3730 -4065 3770 -3995
rect 3730 -4085 3740 -4065
rect 3760 -4085 3770 -4065
rect 3730 -4095 3770 -4085
rect 4330 -4090 4370 -3995
rect 3130 -4120 3170 -4110
rect 4330 -4110 4340 -4090
rect 4360 -4110 4370 -4090
rect 4330 -4120 4370 -4110
rect 4930 -4090 4970 -3995
rect 4930 -4110 4940 -4090
rect 4960 -4110 4970 -4090
rect 4930 -4120 4970 -4110
rect 5530 -4090 5570 -3995
rect 5530 -4110 5540 -4090
rect 5560 -4110 5570 -4090
rect 5530 -4120 5570 -4110
rect 6130 -4090 6170 -3995
rect 6130 -4110 6140 -4090
rect 6160 -4110 6170 -4090
rect 6130 -4120 6170 -4110
rect 6730 -4090 6770 -3995
rect 6730 -4110 6740 -4090
rect 6760 -4110 6770 -4090
rect 6730 -4120 6770 -4110
rect 7330 -4090 7370 -3995
rect 7330 -4110 7340 -4090
rect 7360 -4110 7370 -4090
rect 7330 -4120 7370 -4110
rect 7930 -4090 7970 -3995
rect 7930 -4110 7940 -4090
rect 7960 -4110 7970 -4090
rect 7930 -4120 7970 -4110
<< end >>
