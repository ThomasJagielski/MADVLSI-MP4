magic
tech sky130A
timestamp 1617721049
<< nmos >>
rect -3900 0 -3500 1600
rect -3100 0 -2700 1600
rect -2300 0 -1900 1600
rect -1500 0 -1100 1600
rect -700 0 -300 1600
rect 100 0 500 1600
rect 900 0 1300 1600
rect 1700 0 2100 1600
rect 2500 0 2900 1600
rect 3300 0 3700 1600
rect 4100 0 4500 1600
rect 4900 0 5300 1600
rect 5700 0 6100 1600
rect 6500 0 6900 1600
rect 7300 0 7700 1600
rect 8100 0 8500 1600
rect 8900 0 9300 1600
rect 9700 0 10100 1600
rect 10500 0 10900 1600
rect -3900 -2000 -3500 -400
rect -3100 -2000 -2700 -400
rect -2300 -2000 -1900 -400
rect -1500 -2000 -1100 -400
rect -700 -2000 -300 -400
rect 100 -2000 500 -400
rect 900 -2000 1300 -400
rect 1700 -2000 2100 -400
rect 2500 -2000 2900 -400
rect 3300 -2000 3700 -400
rect 4100 -2000 4500 -400
rect 4900 -2000 5300 -400
rect 5700 -2000 6100 -400
rect 6500 -2000 6900 -400
rect 7300 -2000 7700 -400
rect 8100 -2000 8500 -400
rect 8900 -2000 9300 -400
rect 9700 -2000 10100 -400
rect 10500 -2000 10900 -400
rect -3900 -4000 -3500 -2400
rect -3100 -4000 -2700 -2400
rect -2300 -4000 -1900 -2400
rect -1500 -4000 -1100 -2400
rect -700 -4000 -300 -2400
rect 100 -4000 500 -2400
rect 900 -4000 1300 -2400
rect 1700 -4000 2100 -2400
rect 2500 -4000 2900 -2400
rect 3300 -4000 3700 -2400
rect 4100 -4000 4500 -2400
rect 4900 -4000 5300 -2400
rect 5700 -4000 6100 -2400
rect 6500 -4000 6900 -2400
rect 7300 -4000 7700 -2400
rect 8100 -4000 8500 -2400
rect 8900 -4000 9300 -2400
rect 9700 -4000 10100 -2400
rect 10500 -4000 10900 -2400
<< ndiff >>
rect -4300 1585 -3900 1600
rect -4300 15 -4285 1585
rect -3915 15 -3900 1585
rect -4300 0 -3900 15
rect -3500 1585 -3100 1600
rect -3500 15 -3485 1585
rect -3115 15 -3100 1585
rect -3500 0 -3100 15
rect -2700 1585 -2300 1600
rect -2700 15 -2685 1585
rect -2315 15 -2300 1585
rect -2700 0 -2300 15
rect -1900 1585 -1500 1600
rect -1900 15 -1885 1585
rect -1515 15 -1500 1585
rect -1900 0 -1500 15
rect -1100 1585 -700 1600
rect -1100 15 -1085 1585
rect -715 15 -700 1585
rect -1100 0 -700 15
rect -300 1585 100 1600
rect -300 15 -285 1585
rect 85 15 100 1585
rect -300 0 100 15
rect 500 1585 900 1600
rect 500 15 515 1585
rect 885 15 900 1585
rect 500 0 900 15
rect 1300 1585 1700 1600
rect 1300 15 1315 1585
rect 1685 15 1700 1585
rect 1300 0 1700 15
rect 2100 1585 2500 1600
rect 2100 15 2115 1585
rect 2485 15 2500 1585
rect 2100 0 2500 15
rect 2900 1585 3300 1600
rect 2900 15 2915 1585
rect 3285 15 3300 1585
rect 2900 0 3300 15
rect 3700 1585 4100 1600
rect 3700 15 3715 1585
rect 4085 15 4100 1585
rect 3700 0 4100 15
rect 4500 1585 4900 1600
rect 4500 15 4515 1585
rect 4885 15 4900 1585
rect 4500 0 4900 15
rect 5300 1585 5700 1600
rect 5300 15 5315 1585
rect 5685 15 5700 1585
rect 5300 0 5700 15
rect 6100 1585 6500 1600
rect 6100 15 6115 1585
rect 6485 15 6500 1585
rect 6100 0 6500 15
rect 6900 1585 7300 1600
rect 6900 15 6915 1585
rect 7285 15 7300 1585
rect 6900 0 7300 15
rect 7700 1585 8100 1600
rect 7700 15 7715 1585
rect 8085 15 8100 1585
rect 7700 0 8100 15
rect 8500 1585 8900 1600
rect 8500 15 8515 1585
rect 8885 15 8900 1585
rect 8500 0 8900 15
rect 9300 1585 9700 1600
rect 9300 15 9315 1585
rect 9685 15 9700 1585
rect 9300 0 9700 15
rect 10100 1585 10500 1600
rect 10100 15 10115 1585
rect 10485 15 10500 1585
rect 10100 0 10500 15
rect 10900 1585 11300 1600
rect 10900 15 10915 1585
rect 11285 15 11300 1585
rect 10900 0 11300 15
rect -4300 -415 -3900 -400
rect -4300 -1985 -4285 -415
rect -3915 -1985 -3900 -415
rect -4300 -2000 -3900 -1985
rect -3500 -415 -3100 -400
rect -3500 -1985 -3485 -415
rect -3115 -1985 -3100 -415
rect -3500 -2000 -3100 -1985
rect -2700 -415 -2300 -400
rect -2700 -1985 -2685 -415
rect -2315 -1985 -2300 -415
rect -2700 -2000 -2300 -1985
rect -1900 -415 -1500 -400
rect -1900 -1985 -1885 -415
rect -1515 -1985 -1500 -415
rect -1900 -2000 -1500 -1985
rect -1100 -415 -700 -400
rect -1100 -1985 -1085 -415
rect -715 -1985 -700 -415
rect -1100 -2000 -700 -1985
rect -300 -415 100 -400
rect -300 -1985 -285 -415
rect 85 -1985 100 -415
rect -300 -2000 100 -1985
rect 500 -415 900 -400
rect 500 -1985 515 -415
rect 885 -1985 900 -415
rect 500 -2000 900 -1985
rect 1300 -415 1700 -400
rect 1300 -1985 1315 -415
rect 1685 -1985 1700 -415
rect 1300 -2000 1700 -1985
rect 2100 -415 2500 -400
rect 2100 -1985 2115 -415
rect 2385 -1985 2500 -415
rect 2100 -2000 2500 -1985
rect 2900 -415 3300 -400
rect 2900 -1985 2915 -415
rect 3285 -1985 3300 -415
rect 2900 -2000 3300 -1985
rect 3700 -415 4100 -400
rect 3700 -1985 3715 -415
rect 4085 -1985 4100 -415
rect 3700 -2000 4100 -1985
rect 4500 -415 4900 -400
rect 4500 -1985 4515 -415
rect 4885 -1985 4900 -415
rect 4500 -2000 4900 -1985
rect 5300 -415 5700 -400
rect 5300 -1985 5315 -415
rect 5685 -1985 5700 -415
rect 5300 -2000 5700 -1985
rect 6100 -415 6500 -400
rect 6100 -1985 6115 -415
rect 6485 -1985 6500 -415
rect 6100 -2000 6500 -1985
rect 6900 -415 7300 -400
rect 6900 -1985 6915 -415
rect 7285 -1985 7300 -415
rect 6900 -2000 7300 -1985
rect 7700 -415 8100 -400
rect 7700 -1985 7715 -415
rect 8085 -1985 8100 -415
rect 7700 -2000 8100 -1985
rect 8500 -415 8900 -400
rect 8500 -1985 8515 -415
rect 8885 -1985 8900 -415
rect 8500 -2000 8900 -1985
rect 9300 -415 9700 -400
rect 9300 -1985 9315 -415
rect 9685 -1985 9700 -415
rect 9300 -2000 9700 -1985
rect 10100 -415 10500 -400
rect 10100 -1985 10115 -415
rect 10485 -1985 10500 -415
rect 10100 -2000 10500 -1985
rect 10900 -415 11300 -400
rect 10900 -1985 10915 -415
rect 11285 -1985 11300 -415
rect 10900 -2000 11300 -1985
rect -4300 -2415 -3900 -2400
rect -4300 -3985 -4285 -2415
rect -3915 -3985 -3900 -2415
rect -4300 -4000 -3900 -3985
rect -3500 -2415 -3100 -2400
rect -3500 -3985 -3485 -2415
rect -3115 -3985 -3100 -2415
rect -3500 -4000 -3100 -3985
rect -2700 -2415 -2300 -2400
rect -2700 -3985 -2685 -2415
rect -2315 -3985 -2300 -2415
rect -2700 -4000 -2300 -3985
rect -1900 -2415 -1500 -2400
rect -1900 -3985 -1885 -2415
rect -1515 -3985 -1500 -2415
rect -1900 -4000 -1500 -3985
rect -1100 -2415 -700 -2400
rect -1100 -3985 -1085 -2415
rect -715 -3985 -700 -2415
rect -1100 -4000 -700 -3985
rect -300 -2415 100 -2400
rect -300 -3985 -285 -2415
rect 85 -3985 100 -2415
rect -300 -4000 100 -3985
rect 500 -2415 900 -2400
rect 500 -3985 515 -2415
rect 885 -3985 900 -2415
rect 500 -4000 900 -3985
rect 1300 -2415 1700 -2400
rect 1300 -3985 1315 -2415
rect 1685 -3985 1700 -2415
rect 1300 -4000 1700 -3985
rect 2100 -2415 2500 -2400
rect 2100 -3985 2115 -2415
rect 2385 -3985 2500 -2415
rect 2100 -4000 2500 -3985
rect 2900 -2415 3300 -2400
rect 2900 -3985 2915 -2415
rect 3285 -3985 3300 -2415
rect 2900 -4000 3300 -3985
rect 3700 -2415 4100 -2400
rect 3700 -3985 3715 -2415
rect 4085 -3985 4100 -2415
rect 3700 -4000 4100 -3985
rect 4500 -2415 4900 -2400
rect 4500 -3985 4515 -2415
rect 4885 -3985 4900 -2415
rect 4500 -4000 4900 -3985
rect 5300 -2415 5700 -2400
rect 5300 -3985 5315 -2415
rect 5685 -3985 5700 -2415
rect 5300 -4000 5700 -3985
rect 6100 -2415 6500 -2400
rect 6100 -3985 6115 -2415
rect 6485 -3985 6500 -2415
rect 6100 -4000 6500 -3985
rect 6900 -2415 7300 -2400
rect 6900 -3985 6915 -2415
rect 7285 -3985 7300 -2415
rect 6900 -4000 7300 -3985
rect 7700 -2415 8100 -2400
rect 7700 -3985 7715 -2415
rect 8085 -3985 8100 -2415
rect 7700 -4000 8100 -3985
rect 8500 -2415 8900 -2400
rect 8500 -3985 8515 -2415
rect 8885 -3985 8900 -2415
rect 8500 -4000 8900 -3985
rect 9300 -2415 9700 -2400
rect 9300 -3985 9315 -2415
rect 9685 -3985 9700 -2415
rect 9300 -4000 9700 -3985
rect 10100 -2415 10500 -2400
rect 10100 -3985 10115 -2415
rect 10485 -3985 10500 -2415
rect 10100 -4000 10500 -3985
rect 10900 -2415 11300 -2400
rect 10900 -3985 10915 -2415
rect 11285 -3985 11300 -2415
rect 10900 -4000 11300 -3985
<< ndiffc >>
rect -4285 15 -3915 1585
rect -3485 15 -3115 1585
rect -2685 15 -2315 1585
rect -1885 15 -1515 1585
rect -1085 15 -715 1585
rect -285 15 85 1585
rect 515 15 885 1585
rect 1315 15 1685 1585
rect 2115 15 2485 1585
rect 2915 15 3285 1585
rect 3715 15 4085 1585
rect 4515 15 4885 1585
rect 5315 15 5685 1585
rect 6115 15 6485 1585
rect 6915 15 7285 1585
rect 7715 15 8085 1585
rect 8515 15 8885 1585
rect 9315 15 9685 1585
rect 10115 15 10485 1585
rect 10915 15 11285 1585
rect -4285 -1985 -3915 -415
rect -3485 -1985 -3115 -415
rect -2685 -1985 -2315 -415
rect -1885 -1985 -1515 -415
rect -1085 -1985 -715 -415
rect -285 -1985 85 -415
rect 515 -1985 885 -415
rect 1315 -1985 1685 -415
rect 2115 -1985 2385 -415
rect 2915 -1985 3285 -415
rect 3715 -1985 4085 -415
rect 4515 -1985 4885 -415
rect 5315 -1985 5685 -415
rect 6115 -1985 6485 -415
rect 6915 -1985 7285 -415
rect 7715 -1985 8085 -415
rect 8515 -1985 8885 -415
rect 9315 -1985 9685 -415
rect 10115 -1985 10485 -415
rect 10915 -1985 11285 -415
rect -4285 -3985 -3915 -2415
rect -3485 -3985 -3115 -2415
rect -2685 -3985 -2315 -2415
rect -1885 -3985 -1515 -2415
rect -1085 -3985 -715 -2415
rect -285 -3985 85 -2415
rect 515 -3985 885 -2415
rect 1315 -3985 1685 -2415
rect 2115 -3985 2385 -2415
rect 2915 -3985 3285 -2415
rect 3715 -3985 4085 -2415
rect 4515 -3985 4885 -2415
rect 5315 -3985 5685 -2415
rect 6115 -3985 6485 -2415
rect 6915 -3985 7285 -2415
rect 7715 -3985 8085 -2415
rect 8515 -3985 8885 -2415
rect 9315 -3985 9685 -2415
rect 10115 -3985 10485 -2415
rect 10915 -3985 11285 -2415
<< psubdiff >>
rect -1095 1755 -705 1770
rect -1095 1705 -1080 1755
rect -715 1705 -705 1755
rect -2525 1690 -2475 1705
rect -1095 1690 -705 1705
rect -295 1755 95 1770
rect -295 1705 -280 1755
rect 85 1705 95 1755
rect -295 1690 95 1705
rect 2105 1755 2495 1770
rect 2105 1705 2120 1755
rect 2485 1705 2495 1755
rect 2105 1690 2495 1705
rect 2905 1755 3295 1770
rect 2905 1705 2920 1755
rect 3285 1705 3295 1755
rect 2905 1690 3295 1705
rect 4505 1755 4895 1770
rect 4505 1705 4520 1755
rect 4885 1705 4895 1755
rect 4505 1690 4895 1705
rect 6105 1755 6495 1770
rect 6105 1705 6120 1755
rect 6485 1705 6495 1755
rect 6105 1690 6495 1705
rect 7705 1755 8095 1770
rect 7705 1705 7720 1755
rect 8085 1705 8095 1755
rect 7705 1690 8095 1705
rect 8270 1725 8320 1740
rect 8270 1705 8285 1725
rect 8305 1705 8320 1725
rect 8270 1690 8320 1705
rect -2525 1670 -2510 1690
rect -2490 1670 -2475 1690
rect -2525 1655 -2475 1670
rect -4700 1585 -4300 1600
rect -4700 15 -4685 1585
rect -4315 15 -4300 1585
rect -4700 0 -4300 15
rect 11300 1585 11700 1600
rect 11300 15 11315 1585
rect 11685 15 11700 1585
rect 11300 0 11700 15
rect -2535 -225 -2485 -210
rect -2535 -245 -2520 -225
rect -2500 -245 -2485 -225
rect -2535 -260 -2485 -245
rect -1095 -145 -705 -130
rect -1095 -195 -1080 -145
rect -715 -195 -705 -145
rect -1095 -210 -705 -195
rect 1305 -165 1695 -150
rect 1305 -215 1320 -165
rect 1685 -215 1695 -165
rect 1305 -230 1695 -215
rect 3705 -180 4095 -165
rect 3705 -230 3720 -180
rect 4085 -230 4095 -180
rect 3705 -245 4095 -230
rect 6905 -175 7295 -160
rect 6905 -225 6920 -175
rect 7285 -225 7295 -175
rect 6905 -240 7295 -225
rect 8505 -230 8895 -215
rect 8505 -280 8520 -230
rect 8885 -280 8895 -230
rect 8505 -295 8895 -280
rect -4700 -415 -4300 -400
rect -4700 -1985 -4685 -415
rect -4315 -1985 -4300 -415
rect -4700 -2000 -4300 -1985
rect 11300 -415 11700 -400
rect 11300 -1985 11315 -415
rect 11685 -1985 11700 -415
rect 11300 -2000 11700 -1985
rect -1775 -2335 -1725 -2320
rect -1775 -2355 -1760 -2335
rect -1740 -2355 -1725 -2335
rect -1775 -2370 -1725 -2355
rect -145 -2235 -95 -2220
rect -145 -2255 -130 -2235
rect -110 -2255 -95 -2235
rect -145 -2270 -95 -2255
rect 1305 -2305 1695 -2290
rect 1305 -2355 1320 -2305
rect 1685 -2355 1695 -2305
rect 1305 -2370 1695 -2355
rect 3825 -2330 3875 -2315
rect 3825 -2350 3840 -2330
rect 3860 -2350 3875 -2330
rect 3825 -2365 3875 -2350
rect 6255 -2330 6305 -2315
rect 6255 -2350 6270 -2330
rect 6290 -2350 6305 -2330
rect 6255 -2365 6305 -2350
rect 8625 -2330 8675 -2315
rect 8625 -2350 8640 -2330
rect 8660 -2350 8675 -2330
rect 8625 -2365 8675 -2350
rect -4700 -2415 -4300 -2400
rect -4700 -3985 -4685 -2415
rect -4315 -3985 -4300 -2415
rect -4700 -4000 -4300 -3985
rect 11300 -2415 11700 -2400
rect 11300 -3985 11315 -2415
rect 11685 -3985 11700 -2415
rect 11300 -4000 11700 -3985
rect -975 -4045 -925 -4030
rect -975 -4065 -960 -4045
rect -940 -4065 -925 -4045
rect 1425 -4045 1475 -4030
rect 1425 -4065 1440 -4045
rect 1460 -4065 1475 -4045
rect 3825 -4045 3875 -4030
rect 3825 -4065 3840 -4045
rect 3860 -4065 3875 -4045
rect 6225 -4045 6275 -4030
rect 6225 -4065 6240 -4045
rect 6260 -4065 6275 -4045
rect 8500 -4060 8550 -4055
rect -975 -4080 -925 -4065
rect 1425 -4080 1475 -4065
rect 3825 -4080 3875 -4065
rect 6225 -4080 6275 -4065
rect 8500 -4080 8515 -4060
rect 8535 -4080 8550 -4060
rect -2505 -4100 -2455 -4085
rect 8500 -4095 8550 -4080
rect -2505 -4120 -2490 -4100
rect -2470 -4120 -2455 -4100
rect -2505 -4135 -2455 -4120
<< psubdiffcont >>
rect -1080 1705 -715 1755
rect -280 1705 85 1755
rect 2120 1705 2485 1755
rect 2920 1705 3285 1755
rect 4520 1705 4885 1755
rect 6120 1705 6485 1755
rect 7720 1705 8085 1755
rect 8285 1705 8305 1725
rect -2510 1670 -2490 1690
rect -4685 15 -4315 1585
rect 11315 15 11685 1585
rect -2520 -245 -2500 -225
rect -1080 -195 -715 -145
rect 1320 -215 1685 -165
rect 3720 -230 4085 -180
rect 6920 -225 7285 -175
rect 8520 -280 8885 -230
rect -4685 -1985 -4315 -415
rect 11315 -1985 11685 -415
rect -1760 -2355 -1740 -2335
rect -130 -2255 -110 -2235
rect 1320 -2355 1685 -2305
rect 3840 -2350 3860 -2330
rect 6270 -2350 6290 -2330
rect 8640 -2350 8660 -2330
rect -4685 -3985 -4315 -2415
rect 11315 -3985 11685 -2415
rect -960 -4065 -940 -4045
rect 1440 -4065 1460 -4045
rect 3840 -4065 3860 -4045
rect 6240 -4065 6260 -4045
rect 8515 -4080 8535 -4060
rect -2490 -4120 -2470 -4100
<< poly >>
rect 8915 1705 9300 1715
rect 8915 1685 8925 1705
rect 9290 1685 9300 1705
rect 8915 1655 9300 1685
rect -4295 1645 -2700 1655
rect -4295 1625 -4285 1645
rect -3915 1625 -3485 1645
rect -3115 1625 -2700 1645
rect -4295 1615 -2700 1625
rect -3900 1600 -3500 1615
rect -3100 1600 -2700 1615
rect -2300 1640 9300 1655
rect -2300 1600 -1900 1640
rect -1500 1600 -1100 1640
rect -700 1600 -300 1615
rect 100 1600 500 1640
rect 900 1600 1300 1615
rect 1700 1600 2100 1640
rect 2500 1600 2900 1615
rect 3300 1600 3700 1640
rect 4100 1600 4500 1615
rect 4900 1600 5300 1640
rect 5700 1600 6100 1615
rect 6500 1600 6900 1640
rect 7300 1600 7700 1615
rect 8100 1600 8500 1640
rect 8900 1600 9300 1640
rect 9700 1645 11295 1655
rect 9700 1625 10115 1645
rect 10485 1625 10915 1645
rect 11285 1625 11295 1645
rect 9700 1615 11295 1625
rect 9700 1600 10100 1615
rect 10500 1600 10900 1615
rect -3900 -15 -3500 0
rect -3100 -15 -2700 0
rect -2300 -305 -1900 0
rect -1500 -305 -1100 0
rect -700 -15 -300 0
rect -470 -25 -430 -15
rect -470 -45 -460 -25
rect -440 -45 -430 -25
rect -470 -55 -430 -45
rect 100 -305 500 0
rect 900 -15 1300 0
rect 1130 -25 1170 -15
rect 1130 -45 1140 -25
rect 1160 -45 1170 -25
rect 1130 -55 1170 -45
rect 765 -305 1335 -260
rect 1700 -305 2100 0
rect 2500 -15 2900 0
rect 2630 -25 2670 -15
rect 2630 -45 2640 -25
rect 2660 -45 2670 -25
rect 2630 -55 2670 -45
rect 3300 -305 3700 0
rect 4100 -15 4500 0
rect 4900 -15 5300 0
rect 5700 -15 6100 0
rect 4230 -25 4270 -15
rect 4230 -45 4240 -25
rect 4260 -45 4270 -25
rect 4230 -55 4270 -45
rect 5830 -25 5870 -15
rect 5830 -45 5840 -25
rect 5860 -45 5870 -25
rect 5830 -55 5870 -45
rect 4875 -305 5325 -265
rect 6500 -305 6900 0
rect 7300 -15 7700 0
rect 7430 -25 7470 -15
rect 7430 -45 7440 -25
rect 7460 -45 7470 -25
rect 7430 -55 7470 -45
rect 8100 -305 8500 0
rect 8900 -15 9300 0
rect 9700 -15 10100 0
rect 10500 -15 10900 0
rect -2300 -345 905 -305
rect 1295 -345 4915 -305
rect 5285 -345 8500 -305
rect -4295 -355 -2700 -345
rect -4295 -375 -4285 -355
rect -3915 -375 -3485 -355
rect -3115 -375 -2700 -355
rect -4295 -385 -2700 -375
rect -3900 -400 -3500 -385
rect -3100 -400 -2700 -385
rect -2300 -400 -1900 -345
rect -1500 -400 -1100 -345
rect -700 -400 -300 -345
rect 100 -400 500 -345
rect 1130 -355 1170 -345
rect 1130 -375 1140 -355
rect 1160 -375 1170 -355
rect 1130 -385 1170 -375
rect 900 -400 1300 -385
rect 1700 -400 2100 -345
rect 2500 -400 2900 -345
rect 3300 -400 3700 -345
rect 4100 -400 4500 -345
rect 5030 -355 5070 -345
rect 5030 -375 5040 -355
rect 5060 -375 5070 -355
rect 5030 -385 5070 -375
rect 4900 -400 5300 -385
rect 5700 -400 6100 -345
rect 6500 -400 6900 -345
rect 7300 -400 7700 -345
rect 8100 -400 8500 -345
rect 9305 -355 9695 -345
rect 9305 -370 9315 -355
rect 8900 -375 9315 -370
rect 9685 -370 9695 -355
rect 10105 -355 10495 -345
rect 10105 -370 10115 -355
rect 9685 -375 10115 -370
rect 10485 -370 10495 -355
rect 10905 -355 11295 -345
rect 10905 -370 10915 -355
rect 10485 -375 10915 -370
rect 11285 -375 11295 -355
rect 8900 -385 11295 -375
rect 8900 -400 9300 -385
rect 9700 -400 10100 -385
rect 10500 -400 10900 -385
rect -3900 -2015 -3500 -2000
rect -3100 -2015 -2700 -2000
rect -2300 -2015 -1900 -2000
rect -1500 -2015 -1100 -2000
rect -700 -2015 -300 -2000
rect 100 -2015 500 -2000
rect 900 -2015 1300 -2000
rect 1700 -2015 2100 -2000
rect 2500 -2015 2900 -2000
rect 3300 -2015 3700 -2000
rect 4100 -2015 4500 -2000
rect 4900 -2015 5300 -2000
rect 5700 -2015 6100 -2000
rect 6500 -2015 6900 -2000
rect 7300 -2015 7700 -2000
rect 8100 -2015 8500 -2000
rect 8900 -2015 9300 -2000
rect 9700 -2015 10100 -2000
rect 10500 -2015 10900 -2000
rect -1565 -2025 -1525 -2015
rect -1565 -2045 -1555 -2025
rect -1535 -2045 -1525 -2025
rect -1565 -2345 -1525 -2045
rect 2230 -2025 2270 -2015
rect 2230 -2045 2240 -2025
rect 2260 -2045 2270 -2025
rect -1565 -2365 -1555 -2345
rect -1535 -2365 -1525 -2345
rect -1565 -2375 -1525 -2365
rect 2230 -2355 2270 -2045
rect 6125 -2025 6165 -2015
rect 6125 -2045 6135 -2025
rect 6155 -2045 6165 -2025
rect 6125 -2285 6165 -2045
rect 6125 -2305 6135 -2285
rect 6155 -2305 6165 -2285
rect 6125 -2315 6165 -2305
rect 7725 -2025 7765 -2015
rect 7725 -2045 7735 -2025
rect 7755 -2045 7765 -2025
rect 2230 -2375 2240 -2355
rect 2260 -2375 2270 -2355
rect 7725 -2350 7765 -2045
rect 2230 -2385 2270 -2375
rect 7725 -2370 7735 -2350
rect 7755 -2370 7765 -2350
rect 7725 -2380 7765 -2370
rect -3900 -2400 -3500 -2385
rect -3100 -2400 -2700 -2385
rect -2300 -2400 -1900 -2385
rect -1500 -2400 -1100 -2385
rect -700 -2400 -300 -2385
rect 100 -2400 500 -2385
rect 900 -2400 1300 -2385
rect 1700 -2400 2100 -2385
rect 2500 -2400 2900 -2385
rect 3300 -2400 3700 -2385
rect 4100 -2400 4500 -2385
rect 4900 -2400 5300 -2385
rect 5700 -2400 6100 -2385
rect 6500 -2400 6900 -2385
rect 7300 -2400 7700 -2385
rect 8100 -2400 8500 -2385
rect 8900 -2400 9300 -2385
rect 9700 -2400 10100 -2385
rect 10500 -2400 10900 -2385
rect -3900 -4015 -3500 -4000
rect -3100 -4015 -2700 -4000
rect -2300 -4015 -1900 -4000
rect -1500 -4015 -1100 -4000
rect -4295 -4025 -1100 -4015
rect -4295 -4045 -4285 -4025
rect -3915 -4045 -3485 -4025
rect -3115 -4045 -2685 -4025
rect -2315 -4045 -1885 -4025
rect -1515 -4045 -1100 -4025
rect -4295 -4055 -1100 -4045
rect -700 -4035 -300 -4000
rect -700 -4055 -690 -4035
rect -310 -4055 -300 -4035
rect 100 -4025 500 -4000
rect 100 -4045 110 -4025
rect 490 -4045 500 -4025
rect 100 -4055 500 -4045
rect 900 -4035 1300 -4000
rect 900 -4055 910 -4035
rect 1290 -4055 1300 -4035
rect -700 -4065 -300 -4055
rect 900 -4065 1300 -4055
rect 1700 -4035 2100 -4000
rect 1700 -4055 1710 -4035
rect 2090 -4055 2100 -4035
rect 1700 -4065 2100 -4055
rect 2500 -4035 2900 -4000
rect 2500 -4055 2510 -4035
rect 2890 -4055 2900 -4035
rect 2500 -4065 2900 -4055
rect 3300 -4035 3700 -4000
rect 3300 -4055 3310 -4035
rect 3690 -4055 3700 -4035
rect 3300 -4065 3700 -4055
rect 4100 -4035 4500 -4000
rect 4100 -4055 4110 -4035
rect 4490 -4055 4500 -4035
rect 4100 -4065 4500 -4055
rect 4900 -4035 5300 -4000
rect 4900 -4055 4905 -4035
rect 5290 -4055 5300 -4035
rect 4900 -4065 5300 -4055
rect 5700 -4035 6100 -4000
rect 5700 -4055 5710 -4035
rect 6090 -4055 6100 -4035
rect 5700 -4065 6100 -4055
rect 6500 -4035 6900 -4000
rect 6500 -4055 6510 -4035
rect 6890 -4055 6900 -4035
rect 7300 -4015 7700 -4000
rect 8100 -4015 8500 -4000
rect 8900 -4015 9300 -4000
rect 9700 -4015 10100 -4000
rect 10500 -4015 10900 -4000
rect 7300 -4025 11295 -4015
rect 7300 -4045 7715 -4025
rect 8085 -4045 8585 -4025
rect 8885 -4045 9315 -4025
rect 9685 -4045 10115 -4025
rect 10485 -4045 10915 -4025
rect 11285 -4045 11295 -4025
rect 7300 -4055 11295 -4045
rect 6500 -4065 6900 -4055
<< polycont >>
rect 8925 1685 9290 1705
rect -4285 1625 -3915 1645
rect -3485 1625 -3115 1645
rect 10115 1625 10485 1645
rect 10915 1625 11285 1645
rect -460 -45 -440 -25
rect 1140 -45 1160 -25
rect 2640 -45 2660 -25
rect 4240 -45 4260 -25
rect 5840 -45 5860 -25
rect 7440 -45 7460 -25
rect -4285 -375 -3915 -355
rect -3485 -375 -3115 -355
rect 1140 -375 1160 -355
rect 5040 -375 5060 -355
rect 9315 -375 9685 -355
rect 10115 -375 10485 -355
rect 10915 -375 11285 -355
rect -1555 -2045 -1535 -2025
rect 2240 -2045 2260 -2025
rect -1555 -2365 -1535 -2345
rect 6135 -2045 6155 -2025
rect 6135 -2305 6155 -2285
rect 7735 -2045 7755 -2025
rect 2240 -2375 2260 -2355
rect 7735 -2370 7755 -2350
rect -4285 -4045 -3915 -4025
rect -3485 -4045 -3115 -4025
rect -2685 -4045 -2315 -4025
rect -1885 -4045 -1515 -4025
rect -690 -4055 -310 -4035
rect 110 -4045 490 -4025
rect 910 -4055 1290 -4035
rect 1710 -4055 2090 -4035
rect 2510 -4055 2890 -4035
rect 3310 -4055 3690 -4035
rect 4110 -4055 4490 -4035
rect 4905 -4055 5290 -4035
rect 5710 -4055 6090 -4035
rect 6510 -4055 6890 -4035
rect 7715 -4045 8085 -4025
rect 8585 -4045 8885 -4025
rect 9315 -4045 9685 -4025
rect 10115 -4045 10485 -4025
rect 10915 -4045 11285 -4025
<< locali >>
rect -1095 1755 -705 1770
rect -1095 1705 -1080 1755
rect -715 1705 -705 1755
rect -2520 1690 -2480 1700
rect -1095 1690 -705 1705
rect -295 1755 95 1770
rect -295 1705 -280 1755
rect 85 1705 95 1755
rect -295 1690 95 1705
rect 2105 1755 2495 1770
rect 2105 1705 2120 1755
rect 2485 1705 2495 1755
rect 2105 1690 2495 1705
rect 2905 1755 3295 1770
rect 2905 1705 2920 1755
rect 3285 1705 3295 1755
rect 2905 1690 3295 1705
rect 4505 1755 4895 1770
rect 4505 1705 4520 1755
rect 4885 1705 4895 1755
rect 4505 1690 4895 1705
rect 6105 1755 6495 1770
rect 6105 1705 6120 1755
rect 6485 1705 6495 1755
rect 6105 1690 6495 1705
rect 7705 1755 8095 1770
rect 7705 1705 7720 1755
rect 8085 1705 8095 1755
rect 8505 1740 11700 1780
rect 7705 1690 8095 1705
rect 8275 1725 8315 1735
rect 8275 1705 8285 1725
rect 8305 1705 8315 1725
rect 8275 1695 8315 1705
rect -2520 1670 -2510 1690
rect -2490 1670 -2480 1690
rect -2520 1660 -2480 1670
rect -4295 1645 -3905 1655
rect -4295 1625 -4285 1645
rect -3915 1625 -3905 1645
rect -4295 1595 -3905 1625
rect -4695 1585 -3905 1595
rect -4695 15 -4685 1585
rect -4315 15 -4285 1585
rect -3915 15 -3905 1585
rect -4695 5 -3905 15
rect -3495 1645 -3105 1655
rect -3495 1625 -3485 1645
rect -3115 1625 -3105 1645
rect -3495 1585 -3105 1625
rect -3495 15 -3485 1585
rect -3115 15 -3105 1585
rect -3495 5 -3105 15
rect -2695 1585 -2305 1595
rect -2695 15 -2685 1585
rect -2315 15 -2305 1585
rect -2695 -20 -2305 15
rect -1895 1585 -1505 1595
rect -1895 15 -1885 1585
rect -1515 15 -1505 1585
rect -1895 5 -1505 15
rect -1095 1585 -700 1595
rect -1095 15 -1085 1585
rect -715 15 -700 1585
rect -1095 5 -700 15
rect -295 1585 95 1595
rect -295 15 -285 1585
rect 85 15 95 1585
rect -1095 -20 -705 5
rect -2695 -60 -705 -20
rect -470 -25 -430 -15
rect -470 -45 -460 -25
rect -440 -45 -430 -25
rect -295 -40 95 15
rect 505 1585 895 1595
rect 505 15 515 1585
rect 885 15 895 1585
rect 505 5 895 15
rect 1305 1585 1695 1595
rect 1305 15 1315 1585
rect 1685 15 1695 1585
rect 1305 5 1695 15
rect 2105 1585 2495 1595
rect 2105 15 2115 1585
rect 2485 15 2495 1585
rect 1130 -25 1170 -15
rect -470 -55 -430 -45
rect -2530 -225 -2490 -215
rect -2530 -245 -2520 -225
rect -2500 -245 -2490 -225
rect -2530 -255 -2490 -245
rect -4295 -355 -3905 -345
rect -4295 -375 -4285 -355
rect -3915 -375 -3905 -355
rect -4295 -405 -3905 -375
rect -4695 -415 -3905 -405
rect -4695 -1985 -4685 -415
rect -4315 -1985 -4285 -415
rect -3915 -1985 -3905 -415
rect -4695 -1995 -3905 -1985
rect -3495 -355 -3105 -345
rect -3495 -375 -3485 -355
rect -3115 -375 -3105 -355
rect -3495 -415 -3105 -375
rect -3495 -1985 -3485 -415
rect -3115 -1985 -3105 -415
rect -3495 -1995 -3105 -1985
rect -2695 -415 -2305 -405
rect -2695 -1985 -2685 -415
rect -2315 -1985 -2305 -415
rect -2695 -2080 -2305 -1985
rect -1895 -415 -1505 -60
rect -1095 -145 -705 -130
rect -1095 -195 -1080 -145
rect -715 -195 -705 -145
rect -1095 -210 -705 -195
rect -180 -255 -140 -40
rect 1130 -45 1140 -25
rect 1160 -45 1170 -25
rect 1130 -55 1170 -45
rect 1305 -165 1695 -150
rect 1305 -215 1320 -165
rect 1685 -215 1695 -165
rect 1305 -230 1695 -215
rect -1895 -1985 -1885 -415
rect -1515 -1985 -1505 -415
rect -1895 -2015 -1505 -1985
rect -1095 -295 -140 -255
rect -1095 -405 -705 -295
rect 880 -320 1320 -280
rect 2105 -320 2495 15
rect 2905 1585 3295 1595
rect 2905 15 2915 1585
rect 3285 15 3295 1585
rect 2630 -25 2670 -15
rect 2630 -45 2640 -25
rect 2660 -45 2670 -25
rect 2630 -55 2670 -45
rect -295 -360 920 -320
rect 1130 -355 1170 -345
rect -1095 -415 -700 -405
rect -1095 -1985 -1085 -415
rect -715 -1985 -700 -415
rect -1095 -1995 -700 -1985
rect -295 -415 95 -360
rect 1130 -375 1140 -355
rect 1160 -375 1170 -355
rect 1280 -360 2495 -320
rect 1130 -385 1170 -375
rect -295 -1985 -285 -415
rect 85 -1985 95 -415
rect -295 -1995 95 -1985
rect 505 -415 895 -405
rect 505 -1985 515 -415
rect 885 -1985 895 -415
rect -1565 -2025 -1525 -2015
rect -1565 -2045 -1555 -2025
rect -1535 -2045 -1525 -2025
rect -1565 -2055 -1525 -2045
rect -1095 -2080 -705 -1995
rect 505 -2080 895 -1985
rect -2695 -2120 895 -2080
rect 1305 -415 1695 -405
rect 1305 -1985 1315 -415
rect 1685 -1985 1695 -415
rect 1305 -2080 1695 -1985
rect 2105 -415 2495 -360
rect 2105 -1985 2115 -415
rect 2385 -1985 2495 -415
rect 2105 -2015 2495 -1985
rect 2905 -320 3295 15
rect 3705 1585 4095 1595
rect 3705 15 3715 1585
rect 4085 15 4095 1585
rect 3705 5 4095 15
rect 4505 1585 4895 1595
rect 4505 15 4515 1585
rect 4885 15 4895 1585
rect 4230 -25 4270 -15
rect 4230 -45 4240 -25
rect 4260 -45 4270 -25
rect 4230 -55 4270 -45
rect 3705 -180 4095 -165
rect 3705 -230 3720 -180
rect 4085 -230 4095 -180
rect 3705 -245 4095 -230
rect 4505 -260 4895 15
rect 5305 1585 5695 1595
rect 5305 15 5315 1585
rect 5685 15 5695 1585
rect 5305 5 5695 15
rect 6105 1585 6495 1595
rect 6105 15 6115 1585
rect 6485 15 6495 1585
rect 5830 -25 5870 -15
rect 5830 -45 5840 -25
rect 5860 -45 5870 -25
rect 5830 -55 5870 -45
rect 6105 -260 6495 15
rect 6905 1585 7295 1595
rect 6905 15 6915 1585
rect 7285 15 7295 1585
rect 6905 5 7295 15
rect 7705 1585 8095 1595
rect 7705 15 7715 1585
rect 8085 15 8095 1585
rect 7430 -25 7470 -15
rect 7430 -45 7440 -25
rect 7460 -45 7470 -25
rect 7430 -55 7470 -45
rect 7705 -20 8095 15
rect 8505 1585 8895 1740
rect 8915 1705 11700 1715
rect 8915 1685 8925 1705
rect 9290 1685 11700 1705
rect 8915 1675 11700 1685
rect 10105 1645 10495 1655
rect 10105 1625 10115 1645
rect 10485 1625 10495 1645
rect 8505 15 8515 1585
rect 8885 15 8895 1585
rect 8505 5 8895 15
rect 9305 1585 9695 1595
rect 9305 15 9315 1585
rect 9685 15 9695 1585
rect 9305 -20 9695 15
rect 10105 1585 10495 1625
rect 10105 15 10115 1585
rect 10485 15 10495 1585
rect 10105 5 10495 15
rect 10905 1645 11295 1655
rect 10905 1625 10915 1645
rect 11285 1625 11295 1645
rect 10905 1595 11295 1625
rect 10905 1585 11695 1595
rect 10905 15 10915 1585
rect 11285 15 11315 1585
rect 11685 15 11695 1585
rect 10905 5 11695 15
rect 7705 -60 9695 -20
rect 6905 -175 7295 -160
rect 6905 -225 6920 -175
rect 7285 -225 7295 -175
rect 6905 -240 7295 -225
rect 4505 -300 5320 -260
rect 6105 -300 7295 -260
rect 5280 -320 5320 -300
rect 2905 -360 4895 -320
rect 2905 -415 3295 -360
rect 2905 -1985 2915 -415
rect 3285 -1985 3295 -415
rect 2230 -2025 2270 -2015
rect 2230 -2045 2240 -2025
rect 2260 -2045 2270 -2025
rect 2230 -2055 2270 -2045
rect 2905 -2080 3295 -1985
rect 3705 -415 4095 -405
rect 3705 -1985 3715 -415
rect 4085 -1985 4095 -415
rect 3705 -2015 4095 -1985
rect 4505 -415 4895 -360
rect 5030 -355 5070 -345
rect 5030 -375 5040 -355
rect 5060 -375 5070 -355
rect 5280 -360 6495 -320
rect 5030 -385 5070 -375
rect 4505 -1985 4515 -415
rect 4885 -1985 4895 -415
rect 4505 -1995 4895 -1985
rect 5305 -415 5695 -405
rect 5305 -1985 5315 -415
rect 5685 -1985 5695 -415
rect 1305 -2120 3295 -2080
rect -140 -2235 -100 -2225
rect -140 -2255 -130 -2235
rect -110 -2255 -100 -2235
rect -140 -2265 -100 -2255
rect -1770 -2335 -1730 -2325
rect -1770 -2355 -1760 -2335
rect -1740 -2355 -1730 -2335
rect -1770 -2405 -1730 -2355
rect -1565 -2345 95 -2335
rect -1565 -2365 -1555 -2345
rect -1535 -2365 95 -2345
rect -1565 -2375 95 -2365
rect -4695 -2415 -3905 -2405
rect -4695 -3985 -4685 -2415
rect -4315 -3985 -4285 -2415
rect -3915 -3985 -3905 -2415
rect -4695 -3995 -3905 -3985
rect -4295 -4025 -3905 -3995
rect -4295 -4045 -4285 -4025
rect -3915 -4045 -3905 -4025
rect -4295 -4055 -3905 -4045
rect -3495 -2415 -3105 -2405
rect -3495 -3985 -3485 -2415
rect -3115 -3985 -3105 -2415
rect -3495 -4025 -3105 -3985
rect -3495 -4045 -3485 -4025
rect -3115 -4045 -3105 -4025
rect -3495 -4055 -3105 -4045
rect -2695 -2415 -2305 -2405
rect -2695 -3985 -2685 -2415
rect -2315 -3985 -2305 -2415
rect -2695 -4025 -2305 -3985
rect -2695 -4045 -2685 -4025
rect -2315 -4045 -2305 -4025
rect -2695 -4055 -2305 -4045
rect -1895 -2415 -1505 -2405
rect -1895 -3985 -1885 -2415
rect -1515 -3985 -1505 -2415
rect -1895 -4025 -1505 -3985
rect -1095 -2415 -700 -2405
rect -1095 -3985 -1085 -2415
rect -715 -3985 -700 -2415
rect -1095 -3995 -700 -3985
rect -295 -2415 95 -2375
rect -295 -3985 -285 -2415
rect 85 -3985 95 -2415
rect -295 -3995 95 -3985
rect 505 -2415 895 -2120
rect 505 -3985 515 -2415
rect 885 -3985 895 -2415
rect 505 -3995 895 -3985
rect 1305 -2305 1695 -2290
rect 1305 -2355 1320 -2305
rect 1685 -2355 1695 -2305
rect 1305 -2415 1695 -2355
rect 2230 -2355 2270 -2345
rect 2230 -2375 2240 -2355
rect 2260 -2375 2270 -2355
rect 2230 -2385 2270 -2375
rect 1305 -3985 1315 -2415
rect 1685 -3985 1695 -2415
rect 1305 -3995 1695 -3985
rect 2105 -2415 2495 -2385
rect 2105 -3985 2115 -2415
rect 2385 -3985 2495 -2415
rect 2105 -3995 2495 -3985
rect 2905 -2415 3295 -2120
rect 4055 -2275 4095 -2015
rect 5305 -2080 5695 -1985
rect 6105 -415 6495 -360
rect 6105 -1985 6115 -415
rect 6485 -1985 6495 -415
rect 6105 -2015 6495 -1985
rect 6905 -415 7295 -300
rect 6905 -1985 6915 -415
rect 7285 -1985 7295 -415
rect 6125 -2025 6165 -2015
rect 6125 -2045 6135 -2025
rect 6155 -2045 6165 -2025
rect 6125 -2055 6165 -2045
rect 6905 -2080 7295 -1985
rect 7705 -415 8095 -60
rect 8505 -230 8895 -215
rect 8505 -280 8520 -230
rect 8885 -280 8895 -230
rect 8505 -295 8895 -280
rect 9305 -355 9695 -345
rect 9305 -375 9315 -355
rect 9685 -375 9695 -355
rect 7705 -1985 7715 -415
rect 8085 -1985 8095 -415
rect 7705 -2015 8095 -1985
rect 8505 -415 8895 -405
rect 8505 -1985 8515 -415
rect 8885 -1985 8895 -415
rect 7725 -2025 7765 -2015
rect 7725 -2045 7735 -2025
rect 7755 -2045 7765 -2025
rect 7725 -2055 7765 -2045
rect 8505 -2080 8895 -1985
rect 9305 -415 9695 -375
rect 9305 -1985 9315 -415
rect 9685 -1985 9695 -415
rect 9305 -1995 9695 -1985
rect 10105 -355 10495 -345
rect 10105 -375 10115 -355
rect 10485 -375 10495 -355
rect 10105 -415 10495 -375
rect 10105 -1985 10115 -415
rect 10485 -1985 10495 -415
rect 10105 -1995 10495 -1985
rect 10905 -355 11295 -345
rect 10905 -375 10915 -355
rect 11285 -375 11295 -355
rect 10905 -405 11295 -375
rect 10905 -415 11695 -405
rect 10905 -1985 10915 -415
rect 11285 -1985 11315 -415
rect 11685 -1985 11695 -415
rect 10905 -1995 11695 -1985
rect 5305 -2120 8895 -2080
rect 4055 -2285 6165 -2275
rect 4055 -2305 6135 -2285
rect 6155 -2305 6165 -2285
rect 4055 -2315 6165 -2305
rect 3830 -2330 3870 -2320
rect 3830 -2350 3840 -2330
rect 3860 -2350 3870 -2330
rect 3830 -2405 3870 -2350
rect 2905 -3985 2915 -2415
rect 3285 -3985 3295 -2415
rect 2905 -3995 3295 -3985
rect 3705 -2415 4095 -2405
rect 3705 -3985 3715 -2415
rect 4085 -3985 4095 -2415
rect 3705 -3995 4095 -3985
rect 4505 -2415 4895 -2315
rect 6185 -2340 6225 -2120
rect 4505 -3985 4515 -2415
rect 4885 -3985 4895 -2415
rect 4505 -3995 4895 -3985
rect 5305 -2380 6225 -2340
rect 6260 -2330 6300 -2320
rect 6260 -2350 6270 -2330
rect 6290 -2350 6300 -2330
rect 8630 -2330 8670 -2320
rect 5305 -2415 5695 -2380
rect 6260 -2405 6300 -2350
rect 7725 -2350 7765 -2340
rect 7725 -2360 7735 -2350
rect 6905 -2370 7735 -2360
rect 7755 -2370 7765 -2350
rect 6905 -2380 7765 -2370
rect 8630 -2350 8640 -2330
rect 8660 -2350 8670 -2330
rect 5305 -3985 5315 -2415
rect 5685 -3985 5695 -2415
rect 5305 -3995 5695 -3985
rect 6105 -2415 6495 -2405
rect 6105 -3985 6115 -2415
rect 6485 -3985 6495 -2415
rect 6105 -3995 6495 -3985
rect 6905 -2415 7295 -2380
rect 8630 -2405 8670 -2350
rect 6905 -3985 6915 -2415
rect 7285 -3985 7295 -2415
rect 6905 -3995 7295 -3985
rect 7705 -2415 8095 -2405
rect 7705 -3985 7715 -2415
rect 8085 -3985 8095 -2415
rect -1895 -4045 -1885 -4025
rect -1515 -4045 -1505 -4025
rect -1895 -4055 -1505 -4045
rect -970 -4045 -930 -3995
rect 100 -4025 500 -4015
rect -2500 -4100 -2460 -4055
rect -970 -4065 -960 -4045
rect -940 -4065 -930 -4045
rect -700 -4035 -300 -4025
rect -700 -4055 -690 -4035
rect -310 -4055 -300 -4035
rect 100 -4045 110 -4025
rect 490 -4045 500 -4025
rect 100 -4055 500 -4045
rect 900 -4035 1300 -4025
rect 900 -4055 910 -4035
rect 1290 -4055 1300 -4035
rect -700 -4065 -300 -4055
rect 900 -4065 1300 -4055
rect 1430 -4045 1470 -3995
rect 1430 -4065 1440 -4045
rect 1460 -4065 1470 -4045
rect 1700 -4035 2100 -4025
rect 1700 -4055 1710 -4035
rect 2090 -4055 2100 -4035
rect 1700 -4065 2100 -4055
rect 2500 -4035 2900 -4025
rect 2500 -4055 2510 -4035
rect 2890 -4055 2900 -4035
rect 2500 -4065 2900 -4055
rect 3300 -4035 3700 -4025
rect 3300 -4055 3310 -4035
rect 3690 -4055 3700 -4035
rect 3300 -4065 3700 -4055
rect 3830 -4045 3870 -3995
rect 3830 -4065 3840 -4045
rect 3860 -4065 3870 -4045
rect 4100 -4035 4500 -4025
rect 4100 -4055 4110 -4035
rect 4490 -4055 4500 -4035
rect 4100 -4065 4500 -4055
rect 4900 -4035 5300 -4025
rect 4900 -4055 4905 -4035
rect 5290 -4055 5300 -4035
rect 4900 -4065 5300 -4055
rect 5700 -4035 6100 -4025
rect 5700 -4055 5710 -4035
rect 6090 -4055 6100 -4035
rect 5700 -4065 6100 -4055
rect 6230 -4045 6270 -3995
rect 7705 -4025 8095 -3985
rect 6230 -4065 6240 -4045
rect 6260 -4065 6270 -4045
rect 6500 -4035 6900 -4025
rect 6500 -4055 6510 -4035
rect 6890 -4055 6900 -4035
rect 7705 -4045 7715 -4025
rect 8085 -4045 8095 -4025
rect 7705 -4055 8095 -4045
rect 8505 -2415 8895 -2405
rect 8505 -3985 8515 -2415
rect 8885 -3985 8895 -2415
rect 8505 -4015 8895 -3985
rect 6500 -4065 6900 -4055
rect 8505 -4060 8545 -4015
rect 8575 -4025 8895 -4015
rect 8575 -4045 8585 -4025
rect 8885 -4045 8895 -4025
rect 8575 -4055 8895 -4045
rect 9305 -2415 9695 -2405
rect 9305 -3985 9315 -2415
rect 9685 -3985 9695 -2415
rect 9305 -4025 9695 -3985
rect 9305 -4045 9315 -4025
rect 9685 -4045 9695 -4025
rect 9305 -4055 9695 -4045
rect 10105 -2415 10495 -2405
rect 10105 -3985 10115 -2415
rect 10485 -3985 10495 -2415
rect 10105 -4025 10495 -3985
rect 10105 -4045 10115 -4025
rect 10485 -4045 10495 -4025
rect 10105 -4055 10495 -4045
rect 10905 -2415 11695 -2405
rect 10905 -3985 10915 -2415
rect 11285 -3985 11315 -2415
rect 11685 -3985 11695 -2415
rect 10905 -3995 11695 -3985
rect 10905 -4025 11295 -3995
rect 10905 -4045 10915 -4025
rect 11285 -4045 11295 -4025
rect 10905 -4055 11295 -4045
rect -970 -4075 -930 -4065
rect 1430 -4075 1470 -4065
rect 3830 -4075 3870 -4065
rect 6230 -4075 6270 -4065
rect 8505 -4080 8515 -4060
rect 8535 -4080 8545 -4060
rect 8505 -4090 8545 -4080
rect -2500 -4120 -2490 -4100
rect -2470 -4120 -2460 -4100
rect -2500 -4130 -2460 -4120
<< viali >>
rect -1080 1705 -715 1755
rect -280 1705 85 1755
rect 2120 1705 2485 1755
rect 2920 1705 3285 1755
rect 4520 1705 4885 1755
rect 6120 1705 6485 1755
rect 7720 1705 8085 1755
rect 8285 1705 8305 1725
rect -2510 1670 -2490 1690
rect -4685 15 -4315 1585
rect -4285 15 -3915 1585
rect -3485 15 -3115 1585
rect -1885 15 -1515 1585
rect -460 -45 -440 -25
rect 515 15 885 1585
rect 1315 15 1685 1585
rect -2520 -245 -2500 -225
rect -4685 -1985 -4315 -415
rect -4285 -1985 -3915 -415
rect -3485 -1985 -3115 -415
rect -1080 -195 -715 -145
rect 1140 -45 1160 -25
rect 1320 -215 1685 -165
rect 2640 -45 2660 -25
rect 1140 -375 1160 -355
rect 3715 15 4085 1585
rect 4240 -45 4260 -25
rect 3720 -230 4085 -180
rect 5315 15 5685 1585
rect 5840 -45 5860 -25
rect 7440 -45 7460 -25
rect 10115 15 10485 1585
rect 10915 15 11285 1585
rect 11315 15 11685 1585
rect 6920 -225 7285 -175
rect 5040 -375 5060 -355
rect -130 -2255 -110 -2235
rect -4685 -3985 -4315 -2415
rect -4285 -3985 -3915 -2415
rect -3485 -3985 -3115 -2415
rect -2685 -3985 -2315 -2415
rect -1885 -3985 -1515 -2415
rect -1085 -3985 -715 -2415
rect 1320 -2355 1685 -2305
rect 1315 -3985 1685 -2415
rect 8520 -280 8885 -230
rect 9315 -1985 9685 -415
rect 10115 -1985 10485 -415
rect 10915 -1985 11285 -415
rect 11315 -1985 11685 -415
rect 3715 -3985 4085 -2415
rect 6115 -3985 6485 -2415
rect 7715 -3985 8085 -2415
rect 110 -4045 490 -4025
rect 2510 -4055 2890 -4035
rect 4905 -4055 5290 -4035
rect 8515 -3985 8885 -2415
rect 9315 -3985 9685 -2415
rect 10115 -3985 10485 -2415
rect 10915 -3985 11285 -2415
rect 11315 -3985 11685 -2415
<< metal1 >>
rect -4700 1815 11700 3405
rect -2700 1690 -2300 1735
rect -2700 1670 -2510 1690
rect -2490 1670 -2300 1690
rect -4700 1585 -3105 1595
rect -4700 15 -4685 1585
rect -4315 15 -4285 1585
rect -3915 15 -3485 1585
rect -3115 15 -3105 1585
rect -4700 -400 -3105 15
rect -2700 -225 -2300 1670
rect -1895 1585 -1505 1815
rect -1895 15 -1885 1585
rect -1515 15 -1505 1585
rect -1895 5 -1505 15
rect -1095 1755 -705 1770
rect -1095 1705 -1080 1755
rect -715 1705 -705 1755
rect -2700 -245 -2520 -225
rect -2500 -245 -2300 -225
rect -2700 -400 -2300 -245
rect -1095 -145 -705 1705
rect -295 1755 95 1770
rect -295 1705 -280 1755
rect 85 1705 95 1755
rect -1095 -195 -1080 -145
rect -715 -195 -705 -145
rect -1095 -400 -705 -195
rect -470 -25 -430 -15
rect -470 -45 -460 -25
rect -440 -45 -430 -25
rect -470 -400 -430 -45
rect -295 -400 95 1705
rect 505 1585 895 1815
rect 505 15 515 1585
rect 885 15 895 1585
rect 505 5 895 15
rect 1305 1585 1695 1815
rect 2105 1755 2495 1770
rect 2105 1705 2120 1755
rect 2485 1705 2495 1755
rect 2105 1600 2495 1705
rect 2905 1755 3295 1770
rect 2905 1705 2920 1755
rect 3285 1705 3295 1755
rect 2905 1600 3295 1705
rect 1305 15 1315 1585
rect 1685 15 1695 1585
rect 3705 1585 4095 1815
rect 1305 5 1695 15
rect 1130 -25 1170 -15
rect 1130 -45 1140 -25
rect 1160 -45 1170 -25
rect 1130 -355 1170 -45
rect 1130 -375 1140 -355
rect 1160 -375 1170 -355
rect 1130 -400 1170 -375
rect 1305 -165 1695 -150
rect 1305 -215 1320 -165
rect 1685 -215 1695 -165
rect 1305 -400 1695 -215
rect 2105 -400 2495 1565
rect 2630 -25 2670 -15
rect 2630 -45 2640 -25
rect 2660 -45 2670 -25
rect 2630 -400 2670 -45
rect 2905 -320 3295 1570
rect 3705 15 3715 1585
rect 4085 15 4095 1585
rect 3705 5 4095 15
rect 4505 1755 4895 1770
rect 4505 1705 4520 1755
rect 4885 1705 4895 1755
rect 4230 -25 4270 -15
rect 4230 -45 4240 -25
rect 4260 -45 4270 -25
rect 3705 -180 4095 -165
rect 3705 -230 3720 -180
rect 4085 -230 4095 -180
rect 3705 -320 4095 -230
rect 4230 -320 4270 -45
rect 4505 -320 4895 1705
rect 5305 1585 5695 1815
rect 5305 15 5315 1585
rect 5685 15 5695 1585
rect 5305 5 5695 15
rect 6105 1755 6495 1770
rect 6105 1705 6120 1755
rect 6485 1705 6495 1755
rect 2905 -340 4895 -320
rect 2905 -400 3295 -340
rect 3705 -400 4095 -340
rect 4230 -400 4270 -340
rect 4505 -400 4895 -340
rect 5830 -25 5870 -15
rect 5830 -45 5840 -25
rect 5860 -45 5870 -25
rect 5030 -355 5070 -345
rect 5030 -375 5040 -355
rect 5060 -375 5070 -355
rect 5030 -400 5070 -375
rect 5830 -400 5870 -45
rect 6105 -320 6495 1705
rect 6905 5 7295 1815
rect 7705 1755 8505 1770
rect 7705 1705 7720 1755
rect 8085 1725 8505 1755
rect 8085 1705 8285 1725
rect 8305 1705 8505 1725
rect 7430 -25 7470 -15
rect 7430 -45 7440 -25
rect 7460 -45 7470 -25
rect 6085 -340 6495 -320
rect 6105 -400 6495 -340
rect 6905 -175 7295 -160
rect 6905 -225 6920 -175
rect 7285 -225 7295 -175
rect 6905 -400 7295 -225
rect 7430 -400 7470 -45
rect 7705 -215 8505 1705
rect 10105 1585 11695 1595
rect 10105 15 10115 1585
rect 10485 15 10915 1585
rect 11285 15 11315 1585
rect 11685 15 11695 1585
rect 7705 -230 8895 -215
rect 7705 -280 8520 -230
rect 8885 -280 8895 -230
rect 7705 -400 8895 -280
rect 10105 -400 11695 15
rect -4700 -415 11700 -400
rect -4700 -1985 -4685 -415
rect -4315 -1985 -4285 -415
rect -3915 -1985 -3485 -415
rect -3115 -1985 9315 -415
rect 9685 -1985 10115 -415
rect 10485 -1985 10915 -415
rect 11285 -1985 11315 -415
rect 11685 -1985 11700 -415
rect -4700 -2235 11700 -1985
rect -4700 -2255 -130 -2235
rect -110 -2255 11700 -2235
rect -4700 -2305 11700 -2255
rect -4700 -2355 1320 -2305
rect 1685 -2355 11700 -2305
rect -4700 -2415 11700 -2355
rect -4700 -3985 -4685 -2415
rect -4315 -3985 -4285 -2415
rect -3915 -3985 -3485 -2415
rect -3115 -3985 -2685 -2415
rect -2315 -3985 -1885 -2415
rect -1515 -3985 -1085 -2415
rect -715 -3985 1315 -2415
rect 1685 -3985 3715 -2415
rect 4085 -3985 6115 -2415
rect 6485 -3985 7715 -2415
rect 8085 -3985 8515 -2415
rect 8885 -3985 9315 -2415
rect 9685 -3985 10115 -2415
rect 10485 -3985 10915 -2415
rect 11285 -3985 11315 -2415
rect 11685 -3985 11700 -2415
rect -4700 -3995 11700 -3985
rect 100 -4025 500 -3995
rect 100 -4045 110 -4025
rect 490 -4045 500 -4025
rect 100 -4055 500 -4045
rect 2500 -4035 2900 -3995
rect 2500 -4055 2510 -4035
rect 2890 -4055 2900 -4035
rect 2500 -4065 2900 -4055
rect 4900 -4035 5300 -3995
rect 4900 -4055 4905 -4035
rect 5290 -4055 5300 -4035
rect 4900 -4065 5300 -4055
<< labels >>
rlabel locali 11700 1695 11700 1695 3 Vg
rlabel poly 6650 -4065 6650 -4065 5 b6
rlabel poly 5850 -4065 5850 -4065 5 b5
rlabel poly 4245 -4065 4245 -4065 5 b4
rlabel poly 3450 -4065 3450 -4065 5 b3
rlabel poly 1850 -4065 1850 -4065 5 b2
rlabel poly 1150 -4065 1150 -4065 5 b1
rlabel metal1 -4700 -2215 -4700 -2215 7 GND
rlabel metal1 -4700 2575 -4700 2575 7 VDD
rlabel poly -445 -4065 -445 -4065 5 b0
<< end >>
