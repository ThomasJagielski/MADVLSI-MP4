magic
tech sky130A
timestamp 1617734396
<< nwell >>
rect 7125 1060 7515 1120
<< nmos >>
rect 3530 -6525 3930 -6520
rect 4330 -6525 4730 -6520
rect 5930 -6525 6330 -6520
rect 6730 -6525 7130 -6520
rect 8330 -6525 8730 -6520
rect 9130 -6525 9530 -6520
<< ndiffc >>
rect -14925 -5245 -14905 -5175
rect -13325 -5245 -13305 -5175
rect -12525 -5245 -12505 -5175
rect -10925 -5245 -10905 -5175
rect -10125 -5245 -10105 -5175
rect -8525 -5245 -8505 -5175
rect -7725 -5245 -7705 -5175
<< poly >>
rect -16775 1190 -16370 1225
rect -16775 1170 -16585 1190
rect -16565 1170 -16370 1190
rect -16775 1145 -16370 1170
rect 7125 1105 7515 1115
rect 7125 1085 7135 1105
rect 7505 1085 7515 1105
rect 7125 925 7515 1085
rect 7125 905 7135 925
rect 7505 905 7515 925
rect 7125 895 7515 905
rect 330 -820 735 -790
rect 330 -840 530 -820
rect 550 -840 735 -820
rect 330 -870 735 -840
rect -15645 -5390 -15605 -5380
rect -15645 -5410 -15635 -5390
rect -15615 -5410 -15605 -5390
rect -15645 -5420 -15605 -5410
rect -14145 -5390 -14105 -5380
rect -14145 -5410 -14135 -5390
rect -14115 -5410 -14105 -5390
rect -14145 -5420 -14105 -5410
rect -13145 -5390 -13105 -5380
rect -13145 -5410 -13135 -5390
rect -13115 -5410 -13105 -5390
rect -13145 -5420 -13105 -5410
rect -11490 -5390 -11450 -5380
rect -11490 -5410 -11480 -5390
rect -11460 -5410 -11450 -5390
rect -11490 -5420 -11450 -5410
rect -10645 -5390 -10605 -5380
rect -10645 -5410 -10635 -5390
rect -10615 -5410 -10605 -5390
rect -10645 -5420 -10605 -5410
rect -9145 -5390 -9105 -5380
rect -9145 -5410 -9135 -5390
rect -9115 -5410 -9105 -5390
rect -9145 -5420 -9105 -5410
rect -8395 -5390 -8355 -5380
rect -8395 -5410 -8385 -5390
rect -8365 -5410 -8355 -5390
rect -8395 -5420 -8355 -5410
rect -15620 -5665 -15605 -5420
rect -14120 -5665 -14105 -5420
rect -13120 -5665 -13105 -5420
rect -11465 -5665 -11450 -5420
rect -10620 -5665 -10605 -5420
rect -9120 -5665 -9105 -5420
rect -8370 -5665 -8355 -5420
rect -15645 -5675 -15605 -5665
rect -15645 -5695 -15635 -5675
rect -15615 -5695 -15605 -5675
rect -15645 -5705 -15605 -5695
rect -14145 -5675 -14105 -5665
rect -14145 -5695 -14135 -5675
rect -14115 -5695 -14105 -5675
rect -14145 -5705 -14105 -5695
rect -13145 -5675 -13105 -5665
rect -13145 -5695 -13135 -5675
rect -13115 -5695 -13105 -5675
rect -13145 -5705 -13105 -5695
rect -11490 -5675 -11450 -5665
rect -11490 -5695 -11480 -5675
rect -11460 -5695 -11450 -5675
rect -11490 -5705 -11450 -5695
rect -10645 -5675 -10605 -5665
rect -10645 -5695 -10635 -5675
rect -10615 -5695 -10605 -5675
rect -10645 -5705 -10605 -5695
rect -9145 -5675 -9105 -5665
rect -9145 -5695 -9135 -5675
rect -9115 -5695 -9105 -5675
rect -9145 -5705 -9105 -5695
rect -8395 -5675 -8355 -5665
rect -8395 -5695 -8385 -5675
rect -8365 -5695 -8355 -5675
rect -8395 -5705 -8355 -5695
rect 3530 -6560 3930 -6525
rect 3530 -6580 3540 -6560
rect 3920 -6580 3930 -6560
rect 3530 -6590 3930 -6580
rect 4330 -6560 4730 -6525
rect 4330 -6580 4340 -6560
rect 4720 -6580 4730 -6560
rect 4330 -6590 4730 -6580
rect 5930 -6560 6330 -6525
rect 5930 -6580 5940 -6560
rect 6320 -6580 6330 -6560
rect 5930 -6590 6330 -6580
rect 6730 -6560 7130 -6525
rect 6730 -6580 6740 -6560
rect 7120 -6580 7130 -6560
rect 6730 -6590 7130 -6580
rect 8330 -6560 8730 -6525
rect 8330 -6580 8340 -6560
rect 8720 -6580 8730 -6560
rect 8330 -6590 8730 -6580
rect 9130 -6560 9530 -6525
rect 9130 -6580 9140 -6560
rect 9520 -6580 9530 -6560
rect 9130 -6590 9530 -6580
<< polycont >>
rect -16585 1170 -16565 1190
rect 7135 1085 7505 1105
rect 7135 905 7505 925
rect 530 -840 550 -820
rect -15635 -5410 -15615 -5390
rect -14135 -5410 -14115 -5390
rect -13135 -5410 -13115 -5390
rect -11480 -5410 -11460 -5390
rect -10635 -5410 -10615 -5390
rect -9135 -5410 -9115 -5390
rect -8385 -5410 -8365 -5390
rect -15635 -5695 -15615 -5675
rect -14135 -5695 -14115 -5675
rect -13135 -5695 -13115 -5675
rect -11480 -5695 -11460 -5675
rect -10635 -5695 -10615 -5675
rect -9135 -5695 -9115 -5675
rect -8385 -5695 -8365 -5675
rect 3540 -6580 3920 -6560
rect 4340 -6580 4720 -6560
rect 5940 -6580 6320 -6560
rect 6740 -6580 7120 -6560
rect 8340 -6580 8720 -6560
rect 9140 -6580 9520 -6560
<< locali >>
rect 11515 2930 14320 2960
rect -19520 1330 -16540 1425
rect -22475 -455 -22200 -355
rect -31270 -2790 -30890 -2395
rect -19520 -2660 -19355 1330
rect -16610 1190 -16540 1330
rect -2775 1230 -2125 1270
rect -16610 1170 -16585 1190
rect -16565 1170 -16540 1190
rect -16610 1160 -16540 1170
rect -2775 1165 -2340 1205
rect -2380 -535 -2340 1165
rect -2165 1040 -2125 1230
rect 7125 1105 7515 1180
rect 7125 1085 7135 1105
rect 7505 1085 7515 1105
rect 7125 1075 7515 1085
rect -2165 1020 -2100 1040
rect 9545 1010 9915 1175
rect 9545 960 11525 1010
rect 6325 850 6715 940
rect 7125 925 7515 935
rect 7125 905 7135 925
rect 7505 905 7515 925
rect 7125 895 7515 905
rect 6325 720 9925 850
rect -2380 -575 560 -535
rect 520 -820 560 -575
rect 520 -840 530 -820
rect 550 -840 560 -820
rect 520 -850 560 -840
rect 9535 -930 9925 720
rect 11135 -745 11525 960
rect -19825 -2760 -19355 -2660
rect -22475 -2975 -22110 -2875
rect -13380 -4540 -13360 -4535
rect -15625 -4790 -15250 -4770
rect -44475 -5070 -44405 -4970
rect -15625 -5380 -15605 -4790
rect -15000 -4835 -14960 -4575
rect -14125 -4790 -13675 -4770
rect -15645 -5390 -15605 -5380
rect -15645 -5410 -15635 -5390
rect -15615 -5410 -15605 -5390
rect -15645 -5420 -15605 -5410
rect -15370 -5295 -15185 -5275
rect -15370 -5490 -15345 -5295
rect -14125 -5380 -14105 -4790
rect -13400 -4835 -13360 -4540
rect -13125 -4790 -12840 -4770
rect -14145 -5390 -14105 -5380
rect -14145 -5410 -14135 -5390
rect -14115 -5410 -14105 -5390
rect -14145 -5420 -14105 -5410
rect -13770 -5295 -13685 -5275
rect -13770 -5490 -13745 -5295
rect -13125 -5380 -13105 -4790
rect -12600 -4835 -12560 -4535
rect -11470 -4790 -11215 -4770
rect -13145 -5390 -13105 -5380
rect -13145 -5410 -13135 -5390
rect -13115 -5410 -13105 -5390
rect -13145 -5420 -13105 -5410
rect -12970 -5295 -12885 -5275
rect -12970 -5490 -12945 -5295
rect -11470 -5380 -11450 -4790
rect -11000 -4835 -10960 -4560
rect -10625 -4785 -10400 -4770
rect -10625 -4790 -10425 -4785
rect -11490 -5390 -11450 -5380
rect -11490 -5410 -11480 -5390
rect -11460 -5410 -11450 -5390
rect -11490 -5420 -11450 -5410
rect -11370 -5295 -11285 -5275
rect -11370 -5490 -11345 -5295
rect -10625 -5380 -10605 -4790
rect -10200 -4835 -10160 -4570
rect -9125 -4790 -8860 -4770
rect -10645 -5390 -10605 -5380
rect -10645 -5410 -10635 -5390
rect -10615 -5410 -10605 -5390
rect -10645 -5420 -10605 -5410
rect -10570 -5295 -10485 -5275
rect -10570 -5490 -10545 -5295
rect -9125 -5380 -9105 -4790
rect -8600 -4835 -8560 -4570
rect -8375 -4790 -8050 -4770
rect -9145 -5390 -9105 -5380
rect -9145 -5410 -9135 -5390
rect -9115 -5410 -9105 -5390
rect -9145 -5420 -9105 -5410
rect -8970 -5295 -8885 -5275
rect -8970 -5490 -8945 -5295
rect -8375 -5380 -8355 -4790
rect -7800 -4835 -7760 -4570
rect -8395 -5390 -8355 -5380
rect -8395 -5410 -8385 -5390
rect -8365 -5410 -8355 -5390
rect -8395 -5420 -8355 -5410
rect -8170 -5295 -8085 -5275
rect -8170 -5490 -8145 -5295
rect -19380 -5590 -2710 -5490
rect -19380 -7155 -19270 -5590
rect -19820 -7255 -19270 -7155
rect -15645 -5675 -15605 -5665
rect -15645 -5695 -15635 -5675
rect -15615 -5695 -15605 -5675
rect -15645 -8120 -15605 -5695
rect -14145 -5675 -14105 -5665
rect -14145 -5695 -14135 -5675
rect -14115 -5695 -14105 -5675
rect -14145 -8120 -14105 -5695
rect -13145 -5675 -13105 -5665
rect -13145 -5695 -13135 -5675
rect -13115 -5695 -13105 -5675
rect -13145 -8120 -13105 -5695
rect -11490 -5675 -11450 -5665
rect -11490 -5695 -11480 -5675
rect -11460 -5695 -11450 -5675
rect -11490 -8120 -11450 -5695
rect -10645 -5675 -10605 -5665
rect -10645 -5695 -10635 -5675
rect -10615 -5695 -10605 -5675
rect -10645 -8120 -10605 -5695
rect -9145 -5675 -9105 -5665
rect -9145 -5695 -9135 -5675
rect -9115 -5695 -9105 -5675
rect -9145 -8120 -9105 -5695
rect -8395 -5675 -8355 -5665
rect -8395 -5695 -8385 -5675
rect -8365 -5695 -8355 -5675
rect -8395 -8120 -8355 -5695
rect -2810 -6740 -2710 -5590
rect 1930 -6740 2330 -6550
rect 3530 -6560 3930 -6550
rect 3530 -6580 3540 -6560
rect 3920 -6580 3930 -6560
rect 3530 -6590 3930 -6580
rect 4330 -6560 4730 -6550
rect 4330 -6580 4340 -6560
rect 4720 -6580 4730 -6560
rect 4330 -6590 4730 -6580
rect 5930 -6560 6330 -6550
rect 5930 -6580 5940 -6560
rect 6320 -6580 6330 -6560
rect 5930 -6590 6330 -6580
rect 6730 -6560 7130 -6550
rect 6730 -6580 6740 -6560
rect 7120 -6580 7130 -6560
rect 6730 -6590 7130 -6580
rect 8330 -6560 8730 -6550
rect 8330 -6580 8340 -6560
rect 8720 -6580 8730 -6560
rect 8330 -6590 8730 -6580
rect 9130 -6560 9530 -6550
rect 9130 -6580 9140 -6560
rect 9520 -6580 9530 -6560
rect 9130 -6590 9530 -6580
rect -2810 -6840 2330 -6740
<< viali >>
rect -14925 -5245 -14905 -5175
rect -13325 -5245 -13305 -5175
rect -12525 -5245 -12505 -5175
rect -10925 -5245 -10905 -5175
rect -10125 -5245 -10105 -5175
rect -8525 -5245 -8505 -5175
rect -7725 -5245 -7705 -5175
rect 3540 -6580 3920 -6560
rect 4340 -6580 4720 -6560
rect 5940 -6580 6320 -6560
rect 6740 -6580 7120 -6560
rect 8340 -6580 8720 -6560
rect 9140 -6580 9520 -6560
<< metal1 >>
rect -44480 2055 -44220 2895
rect -19820 1940 -18975 2895
rect -11975 1380 -11575 1385
rect -11975 1310 -11970 1380
rect -11580 1310 -11575 1380
rect -11975 1305 -11575 1310
rect -2935 1300 14320 2895
rect -2070 -295 14320 1300
rect -22880 -5105 -22485 -4855
rect -15285 -4945 -7670 -4830
rect -15285 -5015 -11970 -4945
rect -11580 -5015 -7670 -4945
rect -15285 -5020 -7670 -5015
rect -15285 -5175 -14870 -5100
rect -15285 -5245 -14925 -5175
rect -14905 -5245 -14870 -5175
rect -15285 -5455 -14870 -5245
rect -13685 -5175 -13270 -5075
rect -13685 -5245 -13325 -5175
rect -13305 -5245 -13270 -5175
rect -13685 -5455 -13270 -5245
rect -12885 -5175 -12470 -5115
rect -12885 -5245 -12525 -5175
rect -12505 -5245 -12470 -5175
rect -12885 -5455 -12470 -5245
rect -11285 -5175 -10870 -5085
rect -11285 -5245 -10925 -5175
rect -10905 -5245 -10870 -5175
rect -11285 -5455 -10870 -5245
rect -10485 -5175 -10070 -5090
rect -10485 -5245 -10125 -5175
rect -10105 -5245 -10070 -5175
rect -10485 -5455 -10070 -5245
rect -8885 -5175 -8470 -5085
rect -8885 -5245 -8525 -5175
rect -8505 -5245 -8470 -5175
rect -8885 -5455 -8470 -5245
rect -8085 -5175 -7670 -5105
rect -8085 -5245 -7725 -5175
rect -7705 -5245 -7670 -5175
rect -8085 -5455 -7670 -5245
rect -20905 -6560 14330 -5455
rect -20905 -6580 3540 -6560
rect 3920 -6580 4340 -6560
rect 4720 -6580 5940 -6560
rect 6320 -6580 6740 -6560
rect 7120 -6580 8340 -6560
rect 8720 -6580 9140 -6560
rect 9520 -6580 14330 -6560
rect -44485 -8000 -44030 -7285
rect -20905 -8000 14330 -6580
<< via1 >>
rect -11970 1310 -11580 1380
rect -11970 -5015 -11580 -4945
<< metal2 >>
rect -11975 1380 -11575 1385
rect -11975 1310 -11970 1380
rect -11580 1310 -11575 1380
rect -11975 -4945 -11575 1310
rect -11975 -5015 -11970 -4945
rect -11580 -5015 -11575 -4945
rect -11975 -5020 -11575 -5015
use ibias_vg  ibias_vg_0
timestamp 1617552423
transform 1 0 -43680 0 1 300
box -820 -8300 24030 2600
use mux2  mux2_6
timestamp 1616853209
transform 1 0 -8085 0 1 -5275
box 0 -60 415 505
use mux2  mux2_5
timestamp 1616853209
transform 1 0 -8885 0 1 -5275
box 0 -60 415 505
use mux2  mux2_4
timestamp 1616853209
transform 1 0 -10485 0 1 -5275
box 0 -60 415 505
use mux2  mux2_3
timestamp 1616853209
transform 1 0 -11285 0 1 -5275
box 0 -60 415 505
use mux2  mux2_2
timestamp 1616853209
transform 1 0 -12885 0 1 -5275
box 0 -60 415 505
use mux2  mux2_1
timestamp 1616853209
transform 1 0 -13685 0 1 -5275
box 0 -60 415 505
use mux2  mux2_0
timestamp 1616853209
transform 1 0 -15285 0 1 -5275
box 0 -60 415 505
use low-voltage_super-wilson  low-voltage_super-wilson_0
timestamp 1617552636
transform 1 0 -1485 0 1 1175
box -615 -275 15825 1785
use dac_ladder_wilson  dac_ladder_wilson_0
timestamp 1617721049
transform 1 0 2630 0 1 -2525
box -4700 -4135 11700 3405
use dac_ladder  dac_ladder_0
timestamp 1617561611
transform 1 0 -14475 0 1 -510
box -4700 -4135 11700 3405
<< labels >>
rlabel locali -13685 -5285 -13685 -5285 7 A
rlabel locali -12885 -5285 -12885 -5285 7 A
rlabel locali -11285 -5285 -11285 -5285 7 A
rlabel locali -10485 -5285 -10485 -5285 7 A
rlabel locali -8885 -5285 -8885 -5285 7 A
rlabel locali -8085 -5285 -8085 -5285 7 A
rlabel locali 14320 2945 14320 2945 3 Vout
rlabel locali -44475 -5025 -44475 -5025 7 Vr
rlabel metal1 -44480 2490 -44480 2490 7 VP
rlabel locali -15625 -8120 -15625 -8120 5 s0
rlabel locali -14125 -8120 -14125 -8120 5 s1
rlabel locali -13125 -8120 -13125 -8120 5 s2
rlabel locali -11470 -8120 -11470 -8120 5 s3
rlabel locali -10625 -8120 -10625 -8120 5 s4
rlabel locali -9125 -8120 -9125 -8120 5 s5
rlabel locali -8375 -8120 -8375 -8120 5 s6
rlabel metal1 -18345 -8000 -18345 -8000 5 GND
rlabel locali -19435 1425 -19435 1425 1 Vg
rlabel metal1 -19425 2895 -19425 2895 1 VDD
rlabel locali -30890 -2590 -30890 -2590 3 net10
rlabel metal1 -22485 -4985 -22485 -4985 3 net1
rlabel locali -22325 -355 -22325 -355 1 net2
rlabel locali -22300 -2875 -22300 -2875 1 net3
<< end >>
