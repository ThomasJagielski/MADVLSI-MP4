magic
tech sky130A
timestamp 1617552423
<< nwell >>
rect -820 -2550 17220 1760
<< nmos >>
rect 18800 5 19200 1605
rect 19600 5 20000 1605
rect 20400 5 20800 1605
rect 21200 5 21600 1605
rect 22000 5 22400 1605
rect 22800 5 23200 1605
rect 18800 -2395 19200 -795
rect 19600 -2395 20000 -795
rect 20400 -2395 20800 -795
rect 21200 -2395 21600 -795
rect 22000 -2395 22400 -795
rect 22800 -2395 23200 -795
rect 0 -4915 400 -3315
rect 800 -4915 1200 -3315
rect 1600 -4915 2000 -3315
rect 2400 -4915 2800 -3315
rect 3200 -4915 3600 -3315
rect 4000 -4915 4400 -3315
rect 4800 -4915 5200 -3315
rect 5600 -4915 6000 -3315
rect 6400 -4915 6800 -3315
rect 7200 -4915 7600 -3315
rect 8000 -4915 8400 -3315
rect 8800 -4915 9200 -3315
rect 9600 -4915 10000 -3315
rect 10400 -4915 10800 -3315
rect 12000 -4915 12400 -3315
rect 12800 -4915 13200 -3315
rect 13600 -4915 14000 -3315
rect 14400 -4915 14800 -3315
rect 15200 -4915 15600 -3315
rect 16000 -4915 16400 -3315
rect 18800 -4915 19200 -3315
rect 19600 -4915 20000 -3315
rect 20400 -4915 20800 -3315
rect 21200 -4915 21600 -3315
rect 22000 -4915 22400 -3315
rect 22800 -4915 23200 -3315
rect 0 -7315 400 -5715
rect 800 -7315 1200 -5715
rect 1600 -7315 2000 -5715
rect 2400 -7315 2800 -5715
rect 3200 -7315 3600 -5715
rect 4000 -7315 4400 -5715
rect 4800 -7315 5200 -5715
rect 5600 -7315 6000 -5715
rect 6400 -7315 6800 -5715
rect 7200 -7315 7600 -5715
rect 8000 -7315 8400 -5715
rect 8800 -7315 9200 -5715
rect 9600 -7315 10000 -5715
rect 10400 -7315 10800 -5715
rect 12000 -7315 12400 -5715
rect 12800 -7315 13200 -5715
rect 13600 -7315 14000 -5715
rect 14400 -7315 14800 -5715
rect 15200 -7315 15600 -5715
rect 16000 -7315 16400 -5715
rect 18800 -7315 19200 -5715
rect 19600 -7315 20000 -5715
rect 20400 -7315 20800 -5715
rect 21200 -7315 21600 -5715
rect 22000 -7315 22400 -5715
rect 22800 -7315 23200 -5715
<< pmos >>
rect 0 5 400 1605
rect 800 5 1200 1605
rect 1600 5 2000 1605
rect 2400 5 2800 1605
rect 3200 5 3600 1605
rect 4000 5 4400 1605
rect 4800 5 5200 1605
rect 5600 5 6000 1605
rect 6400 5 6800 1605
rect 7200 5 7600 1605
rect 8000 5 8400 1605
rect 8800 5 9200 1605
rect 9600 5 10000 1605
rect 10400 5 10800 1605
rect 12000 5 12400 1605
rect 12800 5 13200 1605
rect 13600 5 14000 1605
rect 14400 5 14800 1605
rect 15200 5 15600 1605
rect 16000 5 16400 1605
rect 0 -2395 400 -795
rect 800 -2395 1200 -795
rect 1600 -2395 2000 -795
rect 2400 -2395 2800 -795
rect 3200 -2395 3600 -795
rect 4000 -2395 4400 -795
rect 4800 -2395 5200 -795
rect 5600 -2395 6000 -795
rect 6400 -2395 6800 -795
rect 7200 -2395 7600 -795
rect 8000 -2395 8400 -795
rect 8800 -2395 9200 -795
rect 9600 -2395 10000 -795
rect 10400 -2395 10800 -795
rect 12000 -2395 12400 -795
rect 12800 -2395 13200 -795
rect 13600 -2395 14000 -795
rect 14400 -2395 14800 -795
rect 15200 -2395 15600 -795
rect 16000 -2395 16400 -795
<< ndiff >>
rect 18400 1585 18800 1605
rect 18400 25 18420 1585
rect 18780 25 18800 1585
rect 18400 5 18800 25
rect 19200 1585 19600 1605
rect 19200 25 19220 1585
rect 19580 25 19600 1585
rect 19200 5 19600 25
rect 20000 1585 20400 1605
rect 20000 25 20020 1585
rect 20380 25 20400 1585
rect 20000 5 20400 25
rect 20800 1585 21200 1605
rect 20800 25 20820 1585
rect 21180 25 21200 1585
rect 20800 5 21200 25
rect 21600 1585 22000 1605
rect 21600 25 21620 1585
rect 21980 25 22000 1585
rect 21600 5 22000 25
rect 22400 1585 22800 1605
rect 22400 25 22420 1585
rect 22780 25 22800 1585
rect 22400 5 22800 25
rect 23200 1585 23600 1605
rect 23200 25 23220 1585
rect 23580 25 23600 1585
rect 23200 5 23600 25
rect 18400 -815 18800 -795
rect 18400 -2375 18420 -815
rect 18780 -2375 18800 -815
rect 18400 -2395 18800 -2375
rect 19200 -815 19600 -795
rect 19200 -2375 19220 -815
rect 19580 -2375 19600 -815
rect 19200 -2395 19600 -2375
rect 20000 -815 20400 -795
rect 20000 -2375 20020 -815
rect 20380 -2375 20400 -815
rect 20000 -2395 20400 -2375
rect 20800 -815 21200 -795
rect 20800 -2375 20820 -815
rect 21180 -2375 21200 -815
rect 20800 -2395 21200 -2375
rect 21600 -815 22000 -795
rect 21600 -2375 21620 -815
rect 21980 -2375 22000 -815
rect 21600 -2395 22000 -2375
rect 22400 -815 22800 -795
rect 22400 -2375 22420 -815
rect 22780 -2375 22800 -815
rect 22400 -2395 22800 -2375
rect 23200 -815 23600 -795
rect 23200 -2375 23220 -815
rect 23580 -2375 23600 -815
rect 23200 -2395 23600 -2375
rect -400 -3335 0 -3315
rect -400 -4895 -380 -3335
rect -20 -4895 0 -3335
rect -400 -4915 0 -4895
rect 400 -3335 800 -3315
rect 400 -4895 420 -3335
rect 780 -4895 800 -3335
rect 400 -4915 800 -4895
rect 1200 -3335 1600 -3315
rect 1200 -4895 1220 -3335
rect 1580 -4895 1600 -3335
rect 1200 -4915 1600 -4895
rect 2000 -3335 2400 -3315
rect 2000 -4895 2020 -3335
rect 2380 -4895 2400 -3335
rect 2000 -4915 2400 -4895
rect 2800 -3335 3200 -3315
rect 2800 -4895 2820 -3335
rect 3180 -4895 3200 -3335
rect 2800 -4915 3200 -4895
rect 3600 -3335 4000 -3315
rect 3600 -4895 3620 -3335
rect 3980 -4895 4000 -3335
rect 3600 -4915 4000 -4895
rect 4400 -3335 4800 -3315
rect 4400 -4895 4420 -3335
rect 4780 -4895 4800 -3335
rect 4400 -4915 4800 -4895
rect 5200 -3335 5600 -3315
rect 5200 -4895 5220 -3335
rect 5580 -4895 5600 -3335
rect 5200 -4915 5600 -4895
rect 6000 -3335 6400 -3315
rect 6000 -4895 6020 -3335
rect 6380 -4895 6400 -3335
rect 6000 -4915 6400 -4895
rect 6800 -3335 7200 -3315
rect 6800 -4895 6820 -3335
rect 7180 -4895 7200 -3335
rect 6800 -4915 7200 -4895
rect 7600 -3335 8000 -3315
rect 7600 -4895 7620 -3335
rect 7980 -4895 8000 -3335
rect 7600 -4915 8000 -4895
rect 8400 -3335 8800 -3315
rect 8400 -4895 8420 -3335
rect 8780 -4895 8800 -3335
rect 8400 -4915 8800 -4895
rect 9200 -3335 9600 -3315
rect 9200 -4895 9220 -3335
rect 9580 -4895 9600 -3335
rect 9200 -4915 9600 -4895
rect 10000 -3335 10400 -3315
rect 10000 -4895 10020 -3335
rect 10380 -4895 10400 -3335
rect 10000 -4915 10400 -4895
rect 10800 -3335 11200 -3315
rect 11600 -3335 12000 -3315
rect 10800 -4895 10820 -3335
rect 11180 -4895 11200 -3335
rect 11600 -4895 11620 -3335
rect 11980 -4895 12000 -3335
rect 10800 -4915 11200 -4895
rect 11600 -4915 12000 -4895
rect 12400 -3335 12800 -3315
rect 12400 -4895 12420 -3335
rect 12780 -4895 12800 -3335
rect 12400 -4915 12800 -4895
rect 13200 -3335 13600 -3315
rect 13200 -4895 13220 -3335
rect 13580 -4895 13600 -3335
rect 13200 -4915 13600 -4895
rect 14000 -3335 14400 -3315
rect 14000 -4895 14020 -3335
rect 14380 -4895 14400 -3335
rect 14000 -4915 14400 -4895
rect 14800 -3335 15200 -3315
rect 14800 -4895 14820 -3335
rect 15180 -4895 15200 -3335
rect 14800 -4915 15200 -4895
rect 15600 -3335 16000 -3315
rect 15600 -4895 15620 -3335
rect 15980 -4895 16000 -3335
rect 15600 -4915 16000 -4895
rect 16400 -3335 16800 -3315
rect 16400 -4895 16420 -3335
rect 16780 -4895 16800 -3335
rect 16400 -4915 16800 -4895
rect 18400 -3335 18800 -3315
rect 18400 -4895 18420 -3335
rect 18780 -4895 18800 -3335
rect 18400 -4915 18800 -4895
rect 19200 -3335 19600 -3315
rect 19200 -4895 19220 -3335
rect 19580 -4895 19600 -3335
rect 19200 -4915 19600 -4895
rect 20000 -3335 20400 -3315
rect 20000 -4895 20020 -3335
rect 20380 -4895 20400 -3335
rect 20000 -4915 20400 -4895
rect 20800 -3335 21200 -3315
rect 20800 -4895 20820 -3335
rect 21180 -4895 21200 -3335
rect 20800 -4915 21200 -4895
rect 21600 -3335 22000 -3315
rect 21600 -4895 21620 -3335
rect 21980 -4895 22000 -3335
rect 21600 -4915 22000 -4895
rect 22400 -3335 22800 -3315
rect 22400 -4895 22420 -3335
rect 22780 -4895 22800 -3335
rect 22400 -4915 22800 -4895
rect 23200 -3335 23600 -3315
rect 23200 -4895 23220 -3335
rect 23580 -4895 23600 -3335
rect 23200 -4915 23600 -4895
rect -400 -5735 0 -5715
rect -400 -7295 -380 -5735
rect -20 -7295 0 -5735
rect -400 -7315 0 -7295
rect 400 -5735 800 -5715
rect 400 -7295 420 -5735
rect 780 -7295 800 -5735
rect 400 -7315 800 -7295
rect 1200 -5735 1600 -5715
rect 1200 -7295 1220 -5735
rect 1580 -7295 1600 -5735
rect 1200 -7315 1600 -7295
rect 2000 -5735 2400 -5715
rect 2000 -7295 2020 -5735
rect 2380 -7295 2400 -5735
rect 2000 -7315 2400 -7295
rect 2800 -5735 3200 -5715
rect 2800 -7295 2820 -5735
rect 3180 -7295 3200 -5735
rect 2800 -7315 3200 -7295
rect 3600 -5735 4000 -5715
rect 3600 -7295 3620 -5735
rect 3980 -7295 4000 -5735
rect 3600 -7315 4000 -7295
rect 4400 -5735 4800 -5715
rect 4400 -7295 4420 -5735
rect 4780 -7295 4800 -5735
rect 4400 -7315 4800 -7295
rect 5200 -5735 5600 -5715
rect 5200 -7295 5220 -5735
rect 5580 -7295 5600 -5735
rect 5200 -7315 5600 -7295
rect 6000 -5735 6400 -5715
rect 6000 -7295 6020 -5735
rect 6380 -7295 6400 -5735
rect 6000 -7315 6400 -7295
rect 6800 -5735 7200 -5715
rect 6800 -7295 6820 -5735
rect 7180 -7295 7200 -5735
rect 6800 -7315 7200 -7295
rect 7600 -5735 8000 -5715
rect 7600 -7295 7620 -5735
rect 7980 -7295 8000 -5735
rect 7600 -7315 8000 -7295
rect 8400 -5735 8800 -5715
rect 8400 -7295 8420 -5735
rect 8780 -7295 8800 -5735
rect 8400 -7315 8800 -7295
rect 9200 -5735 9600 -5715
rect 9200 -7295 9220 -5735
rect 9580 -7295 9600 -5735
rect 9200 -7315 9600 -7295
rect 10000 -5735 10400 -5715
rect 10000 -7295 10020 -5735
rect 10380 -7295 10400 -5735
rect 10000 -7315 10400 -7295
rect 10800 -5735 11200 -5715
rect 11600 -5735 12000 -5715
rect 10800 -7295 10820 -5735
rect 11180 -7295 11200 -5735
rect 11600 -7295 11620 -5735
rect 11980 -7295 12000 -5735
rect 10800 -7315 11200 -7295
rect 11600 -7315 12000 -7295
rect 12400 -5735 12800 -5715
rect 12400 -7295 12420 -5735
rect 12780 -7295 12800 -5735
rect 12400 -7315 12800 -7295
rect 13200 -5735 13600 -5715
rect 13200 -7295 13220 -5735
rect 13580 -7295 13600 -5735
rect 13200 -7315 13600 -7295
rect 14000 -5735 14400 -5715
rect 14000 -7295 14015 -5735
rect 14380 -7295 14400 -5735
rect 14000 -7315 14400 -7295
rect 14800 -5735 15200 -5715
rect 14800 -7295 14820 -5735
rect 15180 -7295 15200 -5735
rect 14800 -7315 15200 -7295
rect 15600 -5735 16000 -5715
rect 15600 -7295 15620 -5735
rect 15980 -7295 16000 -5735
rect 15600 -7315 16000 -7295
rect 16400 -5735 16800 -5715
rect 16400 -7295 16420 -5735
rect 16780 -7295 16800 -5735
rect 16400 -7315 16800 -7295
rect 18400 -5735 18800 -5715
rect 18400 -7300 18420 -5735
rect 18780 -7300 18800 -5735
rect 18400 -7315 18800 -7300
rect 19200 -5735 19600 -5715
rect 19200 -7295 19220 -5735
rect 19580 -7295 19600 -5735
rect 19200 -7315 19600 -7295
rect 20000 -5735 20400 -5715
rect 20000 -7295 20020 -5735
rect 20380 -7295 20400 -5735
rect 20000 -7315 20400 -7295
rect 20800 -5735 21200 -5715
rect 20800 -7295 20820 -5735
rect 21180 -7295 21200 -5735
rect 20800 -7315 21200 -7295
rect 21600 -5735 22000 -5715
rect 21600 -7295 21620 -5735
rect 21980 -7295 22000 -5735
rect 21600 -7315 22000 -7295
rect 22400 -5735 22800 -5715
rect 22400 -7295 22420 -5735
rect 22780 -7295 22800 -5735
rect 22400 -7315 22800 -7295
rect 23200 -5735 23600 -5715
rect 23200 -7295 23220 -5735
rect 23580 -7295 23600 -5735
rect 23200 -7315 23600 -7295
<< pdiff >>
rect -400 1585 0 1605
rect -400 25 -380 1585
rect -20 25 0 1585
rect -400 5 0 25
rect 400 1585 800 1605
rect 400 25 420 1585
rect 780 25 800 1585
rect 400 5 800 25
rect 1200 1585 1600 1605
rect 1200 25 1220 1585
rect 1580 25 1600 1585
rect 1200 5 1600 25
rect 2000 1585 2400 1605
rect 2000 25 2020 1585
rect 2380 25 2400 1585
rect 2000 5 2400 25
rect 2800 1585 3200 1605
rect 2800 25 2820 1585
rect 3180 25 3200 1585
rect 2800 5 3200 25
rect 3600 1585 4000 1605
rect 3600 25 3620 1585
rect 3980 25 4000 1585
rect 3600 5 4000 25
rect 4400 1585 4800 1605
rect 4400 25 4420 1585
rect 4780 25 4800 1585
rect 4400 5 4800 25
rect 5200 1585 5600 1605
rect 5200 25 5220 1585
rect 5580 25 5600 1585
rect 5200 5 5600 25
rect 6000 1585 6400 1605
rect 6000 25 6020 1585
rect 6380 25 6400 1585
rect 6000 5 6400 25
rect 6800 1585 7200 1605
rect 6800 25 6820 1585
rect 7180 25 7200 1585
rect 6800 5 7200 25
rect 7600 1585 8000 1605
rect 7600 25 7620 1585
rect 7980 25 8000 1585
rect 7600 5 8000 25
rect 8400 1585 8800 1605
rect 8400 25 8420 1585
rect 8780 25 8800 1585
rect 8400 5 8800 25
rect 9200 1585 9600 1605
rect 9200 25 9220 1585
rect 9580 25 9600 1585
rect 9200 5 9600 25
rect 10000 1585 10400 1605
rect 10000 25 10020 1585
rect 10380 25 10400 1585
rect 10000 5 10400 25
rect 10800 1585 11200 1605
rect 11600 1585 12000 1605
rect 10800 25 10820 1585
rect 11180 25 11200 1585
rect 11600 25 11620 1585
rect 11980 25 12000 1585
rect 10800 5 11200 25
rect 11600 5 12000 25
rect 12400 1585 12800 1605
rect 12400 25 12420 1585
rect 12780 25 12800 1585
rect 12400 5 12800 25
rect 13200 1585 13600 1605
rect 13200 25 13220 1585
rect 13580 25 13600 1585
rect 13200 5 13600 25
rect 14000 1585 14400 1605
rect 14000 25 14020 1585
rect 14380 25 14400 1585
rect 14000 5 14400 25
rect 14800 1585 15200 1605
rect 14800 25 14820 1585
rect 15180 25 15200 1585
rect 14800 5 15200 25
rect 15600 1585 16000 1605
rect 15600 25 15620 1585
rect 15980 25 16000 1585
rect 15600 5 16000 25
rect 16400 1585 16800 1605
rect 16400 25 16420 1585
rect 16780 25 16800 1585
rect 16400 5 16800 25
rect -400 -815 0 -795
rect -400 -2375 -380 -815
rect -20 -2375 0 -815
rect -400 -2395 0 -2375
rect 400 -815 800 -795
rect 400 -2375 420 -815
rect 780 -2375 800 -815
rect 400 -2395 800 -2375
rect 1200 -815 1600 -795
rect 1200 -2375 1220 -815
rect 1580 -2375 1600 -815
rect 1200 -2395 1600 -2375
rect 2000 -815 2400 -795
rect 2000 -2375 2020 -815
rect 2380 -2375 2400 -815
rect 2000 -2395 2400 -2375
rect 2800 -815 3200 -795
rect 2800 -2375 2820 -815
rect 3180 -2375 3200 -815
rect 2800 -2395 3200 -2375
rect 3600 -815 4000 -795
rect 3600 -2375 3620 -815
rect 3980 -2375 4000 -815
rect 3600 -2395 4000 -2375
rect 4400 -815 4800 -795
rect 4400 -2375 4420 -815
rect 4780 -2375 4800 -815
rect 4400 -2395 4800 -2375
rect 5200 -815 5600 -795
rect 5200 -2375 5220 -815
rect 5580 -2375 5600 -815
rect 5200 -2395 5600 -2375
rect 6000 -815 6400 -795
rect 6000 -2375 6020 -815
rect 6380 -2375 6400 -815
rect 6000 -2395 6400 -2375
rect 6800 -815 7200 -795
rect 6800 -2375 6820 -815
rect 7180 -2375 7200 -815
rect 6800 -2395 7200 -2375
rect 7600 -815 8000 -795
rect 7600 -2375 7620 -815
rect 7980 -2375 8000 -815
rect 7600 -2395 8000 -2375
rect 8400 -815 8800 -795
rect 8400 -2375 8420 -815
rect 8780 -2375 8800 -815
rect 8400 -2395 8800 -2375
rect 9200 -815 9600 -795
rect 9200 -2375 9220 -815
rect 9580 -2375 9600 -815
rect 9200 -2395 9600 -2375
rect 10000 -815 10400 -795
rect 10000 -2375 10020 -815
rect 10380 -2375 10400 -815
rect 10000 -2395 10400 -2375
rect 10800 -815 11200 -795
rect 11600 -815 12000 -795
rect 10800 -2375 10820 -815
rect 11180 -2375 11200 -815
rect 11600 -2375 11620 -815
rect 11980 -2375 12000 -815
rect 10800 -2395 11200 -2375
rect 11600 -2395 12000 -2375
rect 12400 -815 12800 -795
rect 12400 -2375 12420 -815
rect 12780 -2375 12800 -815
rect 12400 -2395 12800 -2375
rect 13200 -815 13600 -795
rect 13200 -2375 13220 -815
rect 13580 -2375 13600 -815
rect 13200 -2395 13600 -2375
rect 14000 -815 14400 -795
rect 14000 -2375 14020 -815
rect 14380 -2375 14400 -815
rect 14000 -2395 14400 -2375
rect 14800 -815 15200 -795
rect 14800 -2375 14820 -815
rect 15180 -2375 15200 -815
rect 14800 -2395 15200 -2375
rect 15600 -815 16000 -795
rect 15600 -2375 15620 -815
rect 15980 -2375 16000 -815
rect 15600 -2395 16000 -2375
rect 16400 -815 16800 -795
rect 16400 -2375 16420 -815
rect 16780 -2375 16800 -815
rect 16400 -2395 16800 -2375
<< ndiffc >>
rect 18420 25 18780 1585
rect 19220 25 19580 1585
rect 20020 25 20380 1585
rect 20820 25 21180 1585
rect 21620 25 21980 1585
rect 22420 25 22780 1585
rect 23220 25 23580 1585
rect 18420 -2375 18780 -815
rect 19220 -2375 19580 -815
rect 20020 -2375 20380 -815
rect 20820 -2375 21180 -815
rect 21620 -2375 21980 -815
rect 22420 -2375 22780 -815
rect 23220 -2375 23580 -815
rect -380 -4895 -20 -3335
rect 420 -4895 780 -3335
rect 1220 -4895 1580 -3335
rect 2020 -4895 2380 -3335
rect 2820 -4895 3180 -3335
rect 3620 -4895 3980 -3335
rect 4420 -4895 4780 -3335
rect 5220 -4895 5580 -3335
rect 6020 -4895 6380 -3335
rect 6820 -4895 7180 -3335
rect 7620 -4895 7980 -3335
rect 8420 -4895 8780 -3335
rect 9220 -4895 9580 -3335
rect 10020 -4895 10380 -3335
rect 10820 -4895 11180 -3335
rect 11620 -4895 11980 -3335
rect 12420 -4895 12780 -3335
rect 13220 -4895 13580 -3335
rect 14020 -4895 14380 -3335
rect 14820 -4895 15180 -3335
rect 15620 -4895 15980 -3335
rect 16420 -4895 16780 -3335
rect 18420 -4895 18780 -3335
rect 19220 -4895 19580 -3335
rect 20020 -4895 20380 -3335
rect 20820 -4895 21180 -3335
rect 21620 -4895 21980 -3335
rect 22420 -4895 22780 -3335
rect 23220 -4895 23580 -3335
rect -380 -7295 -20 -5735
rect 420 -7295 780 -5735
rect 1220 -7295 1580 -5735
rect 2020 -7295 2380 -5735
rect 2820 -7295 3180 -5735
rect 3620 -7295 3980 -5735
rect 4420 -7295 4780 -5735
rect 5220 -7295 5580 -5735
rect 6020 -7295 6380 -5735
rect 6820 -7295 7180 -5735
rect 7620 -7295 7980 -5735
rect 8420 -7295 8780 -5735
rect 9220 -7295 9580 -5735
rect 10020 -7295 10380 -5735
rect 10820 -7295 11180 -5735
rect 11620 -7295 11980 -5735
rect 12420 -7295 12780 -5735
rect 13220 -7295 13580 -5735
rect 14015 -7295 14380 -5735
rect 14820 -7295 15180 -5735
rect 15620 -7295 15980 -5735
rect 16420 -7295 16780 -5735
rect 18420 -7300 18780 -5735
rect 19220 -7295 19580 -5735
rect 20020 -7295 20380 -5735
rect 20820 -7295 21180 -5735
rect 21620 -7295 21980 -5735
rect 22420 -7295 22780 -5735
rect 23220 -7295 23580 -5735
<< pdiffc >>
rect -380 25 -20 1585
rect 420 25 780 1585
rect 1220 25 1580 1585
rect 2020 25 2380 1585
rect 2820 25 3180 1585
rect 3620 25 3980 1585
rect 4420 25 4780 1585
rect 5220 25 5580 1585
rect 6020 25 6380 1585
rect 6820 25 7180 1585
rect 7620 25 7980 1585
rect 8420 25 8780 1585
rect 9220 25 9580 1585
rect 10020 25 10380 1585
rect 10820 25 11180 1585
rect 11620 25 11980 1585
rect 12420 25 12780 1585
rect 13220 25 13580 1585
rect 14020 25 14380 1585
rect 14820 25 15180 1585
rect 15620 25 15980 1585
rect 16420 25 16780 1585
rect -380 -2375 -20 -815
rect 420 -2375 780 -815
rect 1220 -2375 1580 -815
rect 2020 -2375 2380 -815
rect 2820 -2375 3180 -815
rect 3620 -2375 3980 -815
rect 4420 -2375 4780 -815
rect 5220 -2375 5580 -815
rect 6020 -2375 6380 -815
rect 6820 -2375 7180 -815
rect 7620 -2375 7980 -815
rect 8420 -2375 8780 -815
rect 9220 -2375 9580 -815
rect 10020 -2375 10380 -815
rect 10820 -2375 11180 -815
rect 11620 -2375 11980 -815
rect 12420 -2375 12780 -815
rect 13220 -2375 13580 -815
rect 14020 -2375 14380 -815
rect 14820 -2375 15180 -815
rect 15620 -2375 15980 -815
rect 16420 -2375 16780 -815
<< psubdiff >>
rect 20010 1725 20390 1740
rect 20010 1650 20025 1725
rect 20375 1650 20390 1725
rect 20010 1635 20390 1650
rect 21610 1725 21990 1740
rect 21610 1650 21625 1725
rect 21975 1650 21990 1725
rect 21610 1635 21990 1650
rect 18000 1585 18400 1605
rect 18000 25 18020 1585
rect 18380 25 18400 1585
rect 18000 5 18400 25
rect 23600 1585 24000 1605
rect 23600 25 23620 1585
rect 23980 25 24000 1585
rect 23600 5 24000 25
rect 20010 -400 20390 -385
rect 20010 -475 20025 -400
rect 20375 -475 20390 -400
rect 20010 -490 20390 -475
rect 21620 -385 22000 -370
rect 21620 -460 21635 -385
rect 21985 -460 22000 -385
rect 21620 -475 22000 -460
rect 18000 -815 18400 -795
rect 18000 -2375 18020 -815
rect 18380 -2375 18400 -815
rect 18000 -2395 18400 -2375
rect 23600 -815 24000 -795
rect 23600 -2375 23620 -815
rect 23980 -2375 24000 -815
rect 23600 -2395 24000 -2375
rect 20010 -2780 20390 -2765
rect 20010 -2855 20025 -2780
rect 20375 -2855 20390 -2780
rect 20010 -2870 20390 -2855
rect 2010 -3195 2390 -3180
rect 2010 -3270 2025 -3195
rect 2375 -3270 2390 -3195
rect 2010 -3285 2390 -3270
rect 5210 -3195 5590 -3180
rect 5210 -3270 5225 -3195
rect 5575 -3270 5590 -3195
rect 8410 -3195 8790 -3180
rect 5210 -3285 5590 -3270
rect 8410 -3270 8425 -3195
rect 8775 -3270 8790 -3195
rect 8410 -3285 8790 -3270
rect 14010 -3190 14390 -3175
rect 14010 -3265 14025 -3190
rect 14375 -3265 14390 -3190
rect 14010 -3280 14390 -3265
rect 21610 -2765 21990 -2750
rect 21610 -2840 21625 -2765
rect 21975 -2840 21990 -2765
rect 21610 -2855 21990 -2840
rect -800 -3335 -400 -3315
rect -800 -4895 -780 -3335
rect -420 -4895 -400 -3335
rect -800 -4915 -400 -4895
rect 11200 -3335 11600 -3315
rect 11200 -4895 11220 -3335
rect 11580 -4895 11600 -3335
rect 11200 -4915 11600 -4895
rect 16800 -3335 17200 -3315
rect 16800 -4895 16820 -3335
rect 17180 -4895 17200 -3335
rect 16800 -4915 17200 -4895
rect 18000 -3335 18400 -3315
rect 18000 -4895 18020 -3335
rect 18380 -4895 18400 -3335
rect 18000 -4915 18400 -4895
rect 23600 -3335 24000 -3315
rect 23600 -4895 23620 -3335
rect 23980 -4895 24000 -3335
rect 23600 -4915 24000 -4895
rect 1210 -5145 1590 -5130
rect 1210 -5220 1225 -5145
rect 1575 -5220 1590 -5145
rect 1210 -5235 1590 -5220
rect 4410 -5140 4790 -5125
rect 4410 -5490 4425 -5140
rect 4775 -5490 4790 -5140
rect 4410 -5505 4790 -5490
rect 6410 -5140 6790 -5125
rect 6410 -5490 6425 -5140
rect 6775 -5490 6790 -5140
rect 6410 -5505 6790 -5490
rect 8410 -5140 8790 -5125
rect 8410 -5490 8425 -5140
rect 8775 -5490 8790 -5140
rect 8410 -5505 8790 -5490
rect 14010 -5180 14390 -5165
rect 14010 -5530 14025 -5180
rect 14375 -5530 14390 -5180
rect 14010 -5545 14390 -5530
rect 19265 -5095 19645 -5080
rect 19265 -5445 19280 -5095
rect 19630 -5445 19645 -5095
rect 19265 -5460 19645 -5445
rect 22325 -5110 22705 -5095
rect 22325 -5460 22340 -5110
rect 22690 -5460 22705 -5110
rect 22325 -5475 22705 -5460
rect -800 -5735 -400 -5715
rect -800 -7295 -780 -5735
rect -420 -7295 -400 -5735
rect -800 -7315 -400 -7295
rect 11200 -5735 11600 -5715
rect 11200 -7295 11220 -5735
rect 11580 -7295 11600 -5735
rect 11200 -7315 11600 -7295
rect 16800 -5735 17200 -5715
rect 16800 -7295 16820 -5735
rect 17180 -7295 17200 -5735
rect 16800 -7315 17200 -7295
rect 18000 -5735 18400 -5715
rect 18000 -7295 18020 -5735
rect 18380 -7295 18400 -5735
rect 18000 -7315 18400 -7295
rect 23600 -5735 24000 -5715
rect 23600 -7295 23620 -5735
rect 23980 -7295 24000 -5735
rect 23600 -7315 24000 -7295
rect 2010 -7360 2390 -7345
rect 2010 -7435 2025 -7360
rect 2375 -7435 2390 -7360
rect 2010 -7450 2390 -7435
rect 3610 -7360 3990 -7345
rect 3610 -7435 3625 -7360
rect 3975 -7435 3990 -7360
rect 3610 -7450 3990 -7435
rect 6010 -7360 6390 -7345
rect 6010 -7435 6025 -7360
rect 6375 -7435 6390 -7360
rect 8415 -7360 8785 -7345
rect 8415 -7425 8430 -7360
rect 8770 -7425 8785 -7360
rect 6010 -7450 6390 -7435
rect 8415 -7440 8785 -7425
rect 14015 -7360 14385 -7345
rect 14015 -7425 14030 -7360
rect 14370 -7425 14385 -7360
rect 14015 -7440 14385 -7425
rect 20815 -7360 21185 -7345
rect 20815 -7425 20830 -7360
rect 21170 -7425 21185 -7360
rect 20815 -7440 21185 -7425
<< nsubdiff >>
rect 2010 1725 2390 1740
rect 2010 1650 2025 1725
rect 2375 1650 2390 1725
rect 2010 1635 2390 1650
rect 5210 1725 5590 1740
rect 5210 1650 5225 1725
rect 5575 1650 5590 1725
rect 5210 1635 5590 1650
rect 8410 1725 8790 1740
rect 8410 1650 8425 1725
rect 8775 1650 8790 1725
rect 8410 1635 8790 1650
rect 14010 1725 14390 1740
rect 14010 1650 14025 1725
rect 14375 1650 14390 1725
rect 14010 1635 14390 1650
rect -800 1585 -400 1605
rect -800 25 -780 1585
rect -420 25 -400 1585
rect -800 5 -400 25
rect 11200 1585 11600 1605
rect 11200 25 11220 1585
rect 11580 25 11600 1585
rect 11200 5 11600 25
rect 16800 1585 17200 1605
rect 16800 25 16820 1585
rect 17180 25 17200 1585
rect 16800 5 17200 25
rect 3625 -365 4005 -350
rect 1210 -380 1590 -365
rect 1210 -455 1225 -380
rect 1575 -455 1590 -380
rect 3625 -440 3640 -365
rect 3990 -440 4005 -365
rect 3625 -455 4005 -440
rect 5215 -380 5595 -365
rect 5215 -455 5230 -380
rect 5580 -455 5595 -380
rect 1210 -470 1590 -455
rect 5215 -470 5595 -455
rect 8015 -440 8395 -425
rect 8015 -515 8030 -440
rect 8380 -515 8395 -440
rect 8015 -530 8395 -515
rect 14010 -250 14390 -235
rect 14010 -325 14025 -250
rect 14375 -325 14390 -250
rect 14010 -340 14390 -325
rect -800 -815 -400 -795
rect -800 -2375 -780 -815
rect -420 -2375 -400 -815
rect -800 -2395 -400 -2375
rect 11200 -815 11600 -795
rect 11200 -2375 11220 -815
rect 11580 -2375 11600 -815
rect 11200 -2395 11600 -2375
rect 16800 -815 17200 -795
rect 16800 -2375 16820 -815
rect 17180 -2375 17200 -815
rect 16800 -2395 17200 -2375
rect 2010 -2440 2390 -2425
rect 2010 -2515 2025 -2440
rect 2375 -2515 2390 -2440
rect 2010 -2530 2390 -2515
rect 5210 -2440 5590 -2425
rect 5210 -2515 5225 -2440
rect 5575 -2515 5590 -2440
rect 5210 -2530 5590 -2515
rect 8410 -2440 8790 -2425
rect 8410 -2515 8425 -2440
rect 8775 -2515 8790 -2440
rect 8410 -2530 8790 -2515
rect 14010 -2440 14390 -2425
rect 14010 -2515 14025 -2440
rect 14375 -2515 14390 -2440
rect 14010 -2530 14390 -2515
<< psubdiffcont >>
rect 20025 1650 20375 1725
rect 21625 1650 21975 1725
rect 18020 25 18380 1585
rect 23620 25 23980 1585
rect 20025 -475 20375 -400
rect 21635 -460 21985 -385
rect 18020 -2375 18380 -815
rect 23620 -2375 23980 -815
rect 20025 -2855 20375 -2780
rect 2025 -3270 2375 -3195
rect 5225 -3270 5575 -3195
rect 8425 -3270 8775 -3195
rect 14025 -3265 14375 -3190
rect 21625 -2840 21975 -2765
rect -780 -4895 -420 -3335
rect 11220 -4895 11580 -3335
rect 16820 -4895 17180 -3335
rect 18020 -4895 18380 -3335
rect 23620 -4895 23980 -3335
rect 1225 -5220 1575 -5145
rect 4425 -5490 4775 -5140
rect 6425 -5490 6775 -5140
rect 8425 -5490 8775 -5140
rect 14025 -5530 14375 -5180
rect 19280 -5445 19630 -5095
rect 22340 -5460 22690 -5110
rect -780 -7295 -420 -5735
rect 11220 -7295 11580 -5735
rect 16820 -7295 17180 -5735
rect 18020 -7295 18380 -5735
rect 23620 -7295 23980 -5735
rect 2025 -7435 2375 -7360
rect 3625 -7435 3975 -7360
rect 6025 -7435 6375 -7360
rect 8430 -7425 8770 -7360
rect 14030 -7425 14370 -7360
rect 20830 -7425 21170 -7360
<< nsubdiffcont >>
rect 2025 1650 2375 1725
rect 5225 1650 5575 1725
rect 8425 1650 8775 1725
rect 14025 1650 14375 1725
rect -780 25 -420 1585
rect 11220 25 11580 1585
rect 16820 25 17180 1585
rect 1225 -455 1575 -380
rect 3640 -440 3990 -365
rect 5230 -455 5580 -380
rect 8030 -515 8380 -440
rect 14025 -325 14375 -250
rect -780 -2375 -420 -815
rect 11220 -2375 11580 -815
rect 16820 -2375 17180 -815
rect 2025 -2515 2375 -2440
rect 5225 -2515 5575 -2440
rect 8425 -2515 8775 -2440
rect 14025 -2515 14375 -2440
<< poly >>
rect 4000 1885 6800 1886
rect 3610 1875 6800 1885
rect 3610 1795 3620 1875
rect 3980 1795 6800 1875
rect 3610 1786 6800 1795
rect 3610 1785 4400 1786
rect 3200 1710 3600 1720
rect 3200 1630 3220 1710
rect 3580 1630 3600 1710
rect 0 1605 400 1620
rect 800 1605 1200 1620
rect 1600 1605 2000 1620
rect 2400 1605 2800 1620
rect 3200 1605 3600 1630
rect 4000 1605 4400 1785
rect 4800 1605 5200 1786
rect 5600 1605 6000 1786
rect 6400 1605 6800 1786
rect 7200 1710 7600 1720
rect 7200 1630 7220 1710
rect 7580 1630 7600 1710
rect 7200 1605 7600 1630
rect 8000 1605 8400 1620
rect 8800 1605 9200 1925
rect 9600 1605 10000 1620
rect 10400 1605 10800 1620
rect 12000 1605 12400 1620
rect 12800 1605 13200 1620
rect 13600 1605 14000 1620
rect 14400 1605 14800 1620
rect 15200 1605 15600 1620
rect 16000 1605 16400 1620
rect 18800 1605 19200 1620
rect 19600 1605 20000 1620
rect 20400 1605 20800 1620
rect 21200 1605 21600 1620
rect 22000 1605 22400 1620
rect 22800 1605 23200 1620
rect 0 -10 400 5
rect 800 -10 1200 5
rect -390 -20 1200 -10
rect -390 -100 -380 -20
rect -20 -100 420 -20
rect 780 -100 1200 -20
rect -390 -110 1200 -100
rect 1600 -115 2000 5
rect 2400 -115 2800 5
rect 3200 -10 3600 5
rect 4000 -10 4400 5
rect 4800 -10 5200 5
rect 5600 -10 6000 5
rect 6400 -10 6800 5
rect 7200 -10 7600 5
rect 5820 -20 5990 -10
rect 5820 -80 5830 -20
rect 5980 -80 5990 -20
rect 5820 -90 5990 -80
rect 6410 -20 6580 -10
rect 6410 -80 6420 -20
rect 6570 -80 6580 -20
rect 6410 -90 6580 -80
rect 8000 -115 8400 5
rect 8800 -115 9200 5
rect 9600 -10 10000 5
rect 10400 -10 10800 5
rect 12000 -10 12400 5
rect 9600 -20 11190 -10
rect 9600 -100 10020 -20
rect 10380 -100 10820 -20
rect 11180 -100 11190 -20
rect 9600 -110 11190 -100
rect 11610 -20 12400 -10
rect 11610 -100 11620 -20
rect 11980 -100 12400 -20
rect 11610 -110 12400 -100
rect 1600 -125 9200 -115
rect 1600 -205 6820 -125
rect 7180 -205 9200 -125
rect 1600 -215 9200 -205
rect 12800 -655 13200 5
rect 13600 -655 14000 5
rect 14400 -655 14800 5
rect 15200 -655 15600 5
rect 16000 -10 16400 5
rect 18800 -10 19200 5
rect 16000 -20 16790 -10
rect 16000 -100 16420 -20
rect 16780 -100 16790 -20
rect 16000 -110 16790 -100
rect 18410 -20 19200 -10
rect 18410 -100 18420 -20
rect 18780 -100 19200 -20
rect 18410 -110 19200 -100
rect 12410 -665 15600 -655
rect 3200 -690 3600 -680
rect 3200 -770 3220 -690
rect 3580 -770 3600 -690
rect 7200 -690 7600 -680
rect 0 -795 400 -780
rect 800 -795 1200 -780
rect 1600 -795 2000 -780
rect 2400 -795 2800 -780
rect 3200 -795 3600 -770
rect 5820 -710 5990 -700
rect 5820 -770 5830 -710
rect 5980 -770 5990 -710
rect 5820 -780 5990 -770
rect 6410 -710 6580 -700
rect 6410 -770 6420 -710
rect 6570 -770 6580 -710
rect 6410 -780 6580 -770
rect 7200 -770 7220 -690
rect 7580 -770 7600 -690
rect 12410 -745 12420 -665
rect 12780 -745 15600 -665
rect 12410 -755 15600 -745
rect 4000 -795 4400 -780
rect 4800 -795 5200 -780
rect 5600 -795 6000 -780
rect 6400 -795 6800 -780
rect 7200 -795 7600 -770
rect 8000 -795 8400 -780
rect 8800 -795 9200 -780
rect 9600 -795 10000 -780
rect 10400 -795 10800 -780
rect 12000 -795 12400 -780
rect 12800 -795 13200 -755
rect 13600 -795 14000 -755
rect 14400 -795 14800 -755
rect 15200 -795 15600 -755
rect 16000 -795 16400 -780
rect 18800 -795 19200 -780
rect 19600 -795 20000 5
rect 20400 -795 20800 5
rect 21200 -795 21600 5
rect 22000 -795 22400 5
rect 22800 -10 23200 5
rect 22800 -20 23590 -10
rect 22800 -100 23220 -20
rect 23580 -100 23590 -20
rect 22800 -110 23590 -100
rect 22800 -795 23200 -780
rect 0 -2410 400 -2395
rect 800 -2410 1200 -2395
rect -390 -2420 1200 -2410
rect -390 -2500 -380 -2420
rect -20 -2500 420 -2420
rect 780 -2500 1200 -2420
rect -390 -2510 1200 -2500
rect 1600 -2700 2000 -2395
rect 2400 -2700 2800 -2395
rect 3200 -2410 3600 -2395
rect 4000 -2450 4400 -2395
rect 3610 -2460 4400 -2450
rect 3610 -2540 3620 -2460
rect 3980 -2540 4400 -2460
rect 3610 -2550 4400 -2540
rect 4000 -2575 4400 -2550
rect 4800 -2575 5200 -2395
rect 5600 -2575 6000 -2395
rect 6400 -2575 6800 -2395
rect 7200 -2410 7600 -2395
rect 4000 -2675 6800 -2575
rect 8000 -2700 8400 -2395
rect 8800 -2700 9200 -2395
rect 9600 -2410 10000 -2395
rect 10400 -2410 10800 -2395
rect 12000 -2410 12400 -2395
rect 12800 -2410 13200 -2395
rect 13600 -2410 14000 -2395
rect 14400 -2410 14800 -2395
rect 15200 -2410 15600 -2395
rect 16000 -2410 16400 -2395
rect 18800 -2410 19200 -2395
rect 9600 -2420 11190 -2410
rect 9600 -2500 10020 -2420
rect 10380 -2500 10820 -2420
rect 11180 -2500 11190 -2420
rect 9600 -2510 11190 -2500
rect 11610 -2420 12400 -2410
rect 11610 -2500 11620 -2420
rect 11980 -2500 12400 -2420
rect 16000 -2420 16790 -2410
rect 11610 -2510 12400 -2500
rect 16000 -2500 16420 -2420
rect 16780 -2500 16790 -2420
rect 16000 -2510 16790 -2500
rect 18410 -2420 19200 -2410
rect 18410 -2500 18420 -2420
rect 18780 -2500 19200 -2420
rect 18410 -2510 19200 -2500
rect 1600 -2710 9200 -2700
rect 1600 -2790 6820 -2710
rect 7180 -2790 9200 -2710
rect 1600 -2800 9200 -2790
rect 19600 -2970 20000 -2395
rect 19600 -3050 19610 -2970
rect 19990 -3050 20000 -2970
rect 4000 -3190 4790 -3180
rect 4000 -3270 4420 -3190
rect 4780 -3270 4790 -3190
rect 4000 -3280 4790 -3270
rect 0 -3315 400 -3300
rect 800 -3315 1200 -3300
rect 1600 -3315 2000 -3300
rect 2400 -3315 2800 -3300
rect 3200 -3315 3600 -3300
rect 4000 -3315 4400 -3280
rect 7200 -3270 7600 -3260
rect 7200 -3290 7570 -3270
rect 7590 -3290 7600 -3270
rect 4800 -3315 5200 -3300
rect 5600 -3315 6000 -3300
rect 6400 -3315 6800 -3300
rect 7200 -3315 7600 -3290
rect 8000 -3315 8400 -3300
rect 8800 -3315 9200 -3300
rect 9600 -3315 10000 -3300
rect 10400 -3315 10800 -3300
rect 12000 -3315 12400 -3300
rect 12800 -3315 13200 -3300
rect 13600 -3315 14000 -3300
rect 14400 -3315 14800 -3300
rect 15200 -3315 15600 -3300
rect 16000 -3315 16400 -3300
rect 18800 -3315 19200 -3300
rect 19600 -3315 20000 -3050
rect 20400 -2970 20800 -2395
rect 20400 -3050 20410 -2970
rect 20790 -3050 20800 -2970
rect 20400 -3315 20800 -3050
rect 21200 -2970 21600 -2395
rect 21200 -3050 21210 -2970
rect 21590 -3050 21600 -2970
rect 21200 -3315 21600 -3050
rect 22000 -2970 22400 -2395
rect 22800 -2410 23200 -2395
rect 22800 -2420 23590 -2410
rect 22800 -2500 23220 -2420
rect 23580 -2500 23590 -2420
rect 22800 -2510 23590 -2500
rect 22000 -3050 22010 -2970
rect 22390 -3050 22400 -2970
rect 22000 -3315 22400 -3050
rect 22800 -3315 23200 -3300
rect 0 -4930 400 -4915
rect -390 -4940 400 -4930
rect -390 -5020 -380 -4940
rect -20 -5020 400 -4940
rect -390 -5030 400 -5020
rect 800 -4995 1200 -4915
rect 1600 -4995 2000 -4915
rect 2400 -4995 2800 -4915
rect 3200 -4995 3600 -4915
rect 4000 -4930 4400 -4915
rect 4000 -4940 4450 -4930
rect 4000 -4960 4420 -4940
rect 4440 -4960 4450 -4940
rect 4000 -4970 4450 -4960
rect 4800 -4995 5200 -4915
rect 5600 -4995 6000 -4915
rect 800 -5005 6000 -4995
rect 800 -5085 1220 -5005
rect 1580 -5085 2820 -5005
rect 3180 -5085 6000 -5005
rect 6400 -4940 6800 -4915
rect 6400 -5025 6420 -4940
rect 6780 -5025 6800 -4940
rect 6400 -5035 6800 -5025
rect 7200 -4995 7600 -4915
rect 8000 -4995 8400 -4915
rect 8800 -4995 9200 -4915
rect 9600 -4995 10000 -4915
rect 800 -5095 6000 -5085
rect 800 -5535 1200 -5095
rect 1600 -5535 2000 -5095
rect 2400 -5535 2800 -5095
rect 3200 -5535 3600 -5095
rect 4800 -5535 5200 -5095
rect 5600 -5535 6000 -5095
rect 7200 -5095 10000 -4995
rect 10400 -4930 10800 -4915
rect 12000 -4930 12400 -4915
rect 10400 -4940 11190 -4930
rect 10400 -5020 10820 -4940
rect 11180 -5020 11190 -4940
rect 10400 -5030 11190 -5020
rect 11610 -4940 12400 -4930
rect 11610 -5020 11620 -4940
rect 11980 -5020 12400 -4940
rect 11610 -5030 12400 -5020
rect 800 -5545 6000 -5535
rect 800 -5625 1220 -5545
rect 1580 -5625 2820 -5545
rect 3180 -5625 6000 -5545
rect 7200 -5535 7600 -5095
rect 8000 -5535 8400 -5095
rect 8800 -5535 9200 -5095
rect 9600 -5535 10000 -5095
rect 12800 -5535 13200 -4915
rect 800 -5635 6000 -5625
rect 0 -5715 400 -5700
rect 800 -5715 1200 -5635
rect 1600 -5715 2000 -5635
rect 2400 -5715 2800 -5635
rect 3200 -5715 3600 -5635
rect 4000 -5670 4450 -5660
rect 4000 -5690 4420 -5670
rect 4440 -5690 4450 -5670
rect 4000 -5700 4450 -5690
rect 4000 -5715 4400 -5700
rect 4800 -5715 5200 -5635
rect 5600 -5715 6000 -5635
rect 6400 -5605 6800 -5595
rect 6400 -5690 6420 -5605
rect 6780 -5690 6800 -5605
rect 6400 -5715 6800 -5690
rect 7200 -5635 13200 -5535
rect 7200 -5715 7600 -5635
rect 8000 -5715 8400 -5635
rect 8800 -5715 9200 -5635
rect 9600 -5645 10050 -5635
rect 9600 -5665 10020 -5645
rect 10040 -5665 10050 -5645
rect 9600 -5675 10050 -5665
rect 9600 -5715 10000 -5675
rect 10400 -5715 10800 -5700
rect 12000 -5715 12400 -5700
rect 12800 -5715 13200 -5635
rect 13600 -5715 14000 -4915
rect 14400 -5545 14800 -4915
rect 15200 -5545 15600 -4915
rect 16000 -4930 16400 -4915
rect 18800 -4930 19200 -4915
rect 19600 -4930 20000 -4915
rect 20400 -4930 20800 -4915
rect 21200 -4930 21600 -4915
rect 22000 -4930 22400 -4915
rect 22800 -4930 23200 -4915
rect 16000 -4940 16790 -4930
rect 16000 -5020 16420 -4940
rect 16780 -5020 16790 -4940
rect 16000 -5030 16790 -5020
rect 18410 -4940 19200 -4930
rect 18410 -5020 18420 -4940
rect 18780 -5020 19200 -4940
rect 18410 -5030 19200 -5020
rect 22800 -4940 23590 -4930
rect 22800 -5020 23220 -4940
rect 23580 -5020 23590 -4940
rect 22800 -5030 23590 -5020
rect 14395 -5555 21190 -5545
rect 14395 -5635 20820 -5555
rect 21180 -5635 21190 -5555
rect 14395 -5645 21190 -5635
rect 14400 -5715 14800 -5645
rect 15200 -5715 15600 -5645
rect 16000 -5715 16400 -5700
rect 18800 -5715 19200 -5700
rect 19600 -5715 20000 -5700
rect 20400 -5715 20800 -5700
rect 21200 -5715 21600 -5700
rect 22000 -5715 22400 -5700
rect 22800 -5715 23200 -5700
rect 0 -7330 400 -7315
rect 800 -7330 1200 -7315
rect 1600 -7330 2000 -7315
rect 2400 -7330 2800 -7315
rect 3200 -7330 3600 -7315
rect -390 -7340 400 -7330
rect -390 -7420 -380 -7340
rect -20 -7420 400 -7340
rect -390 -7430 400 -7420
rect 4000 -7350 4400 -7315
rect 4800 -7330 5200 -7315
rect 5600 -7330 6000 -7315
rect 6400 -7330 6800 -7315
rect 7200 -7340 7600 -7315
rect 4000 -7360 4790 -7350
rect 4000 -7440 4420 -7360
rect 4780 -7440 4790 -7360
rect 4000 -7450 4790 -7440
rect 7200 -7420 7210 -7340
rect 7590 -7420 7600 -7340
rect 7200 -7430 7600 -7420
rect 8000 -7340 8400 -7315
rect 8000 -7420 8010 -7340
rect 8390 -7420 8400 -7340
rect 8800 -7340 9200 -7315
rect 8000 -7430 8400 -7420
rect 8800 -7420 8810 -7340
rect 9190 -7420 9200 -7340
rect 8800 -7430 9200 -7420
rect 9600 -7340 10000 -7315
rect 9600 -7420 9610 -7340
rect 9990 -7420 10000 -7340
rect 9600 -7430 10000 -7420
rect 10400 -7330 10800 -7315
rect 12000 -7330 12400 -7315
rect 10400 -7340 11190 -7330
rect 10400 -7420 10820 -7340
rect 11180 -7420 11190 -7340
rect 10400 -7430 11190 -7420
rect 11610 -7340 12400 -7330
rect 11610 -7420 11620 -7340
rect 11980 -7420 12400 -7340
rect 11610 -7430 12400 -7420
rect 12800 -7340 13200 -7315
rect 12800 -7420 12810 -7340
rect 13190 -7420 13200 -7340
rect 12800 -7430 13200 -7420
rect 13600 -7340 14000 -7315
rect 14400 -7330 14800 -7315
rect 15200 -7330 15600 -7315
rect 16000 -7330 16400 -7315
rect 18800 -7330 19200 -7315
rect 13600 -7420 13610 -7340
rect 13990 -7420 14000 -7340
rect 16000 -7340 16790 -7330
rect 13600 -7430 14000 -7420
rect 16000 -7420 16420 -7340
rect 16780 -7420 16790 -7340
rect 16000 -7430 16790 -7420
rect 18410 -7340 19200 -7330
rect 18410 -7420 18420 -7340
rect 18780 -7420 19200 -7340
rect 18410 -7430 19200 -7420
rect 19600 -7340 20000 -7315
rect 19600 -7420 19610 -7340
rect 19990 -7420 20000 -7340
rect 19600 -7430 20000 -7420
rect 20400 -7340 20800 -7315
rect 20400 -7420 20410 -7340
rect 20790 -7420 20800 -7340
rect 21200 -7340 21600 -7315
rect 20400 -7430 20800 -7420
rect 21200 -7420 21210 -7340
rect 21590 -7420 21600 -7340
rect 21200 -7430 21600 -7420
rect 22000 -7340 22400 -7315
rect 22000 -7420 22010 -7340
rect 22390 -7420 22400 -7340
rect 22000 -7430 22400 -7420
rect 22800 -7330 23200 -7315
rect 22800 -7340 23590 -7330
rect 22800 -7420 23220 -7340
rect 23580 -7420 23590 -7340
rect 22800 -7430 23590 -7420
<< polycont >>
rect 3620 1795 3980 1875
rect 3220 1630 3580 1710
rect 7220 1630 7580 1710
rect -380 -100 -20 -20
rect 420 -100 780 -20
rect 5830 -80 5980 -20
rect 6420 -80 6570 -20
rect 10020 -100 10380 -20
rect 10820 -100 11180 -20
rect 11620 -100 11980 -20
rect 6820 -205 7180 -125
rect 16420 -100 16780 -20
rect 18420 -100 18780 -20
rect 3220 -770 3580 -690
rect 5830 -770 5980 -710
rect 6420 -770 6570 -710
rect 7220 -770 7580 -690
rect 12420 -745 12780 -665
rect 23220 -100 23580 -20
rect -380 -2500 -20 -2420
rect 420 -2500 780 -2420
rect 3620 -2540 3980 -2460
rect 10020 -2500 10380 -2420
rect 10820 -2500 11180 -2420
rect 11620 -2500 11980 -2420
rect 16420 -2500 16780 -2420
rect 18420 -2500 18780 -2420
rect 6820 -2790 7180 -2710
rect 19610 -3050 19990 -2970
rect 4420 -3270 4780 -3190
rect 7570 -3290 7590 -3270
rect 20410 -3050 20790 -2970
rect 21210 -3050 21590 -2970
rect 23220 -2500 23580 -2420
rect 22010 -3050 22390 -2970
rect -380 -5020 -20 -4940
rect 4420 -4960 4440 -4940
rect 1220 -5085 1580 -5005
rect 2820 -5085 3180 -5005
rect 6420 -5025 6780 -4940
rect 10820 -5020 11180 -4940
rect 11620 -5020 11980 -4940
rect 1220 -5625 1580 -5545
rect 2820 -5625 3180 -5545
rect 4420 -5690 4440 -5670
rect 6420 -5690 6780 -5605
rect 10020 -5665 10040 -5645
rect 16420 -5020 16780 -4940
rect 18420 -5020 18780 -4940
rect 23220 -5020 23580 -4940
rect 20820 -5635 21180 -5555
rect -380 -7420 -20 -7340
rect 4420 -7440 4780 -7360
rect 7210 -7420 7590 -7340
rect 8010 -7420 8390 -7340
rect 8810 -7420 9190 -7340
rect 9610 -7420 9990 -7340
rect 10820 -7420 11180 -7340
rect 11620 -7420 11980 -7340
rect 12810 -7420 13190 -7340
rect 13610 -7420 13990 -7340
rect 16420 -7420 16780 -7340
rect 18420 -7420 18780 -7340
rect 19610 -7420 19990 -7340
rect 20410 -7420 20790 -7340
rect 21210 -7420 21590 -7340
rect 22010 -7420 22390 -7340
rect 23220 -7420 23580 -7340
<< locali >>
rect 3610 1875 3990 1885
rect 3610 1795 3620 1875
rect 3980 1795 3990 1875
rect 2015 1725 2385 1735
rect 2015 1650 2025 1725
rect 2375 1650 2385 1725
rect 2015 1640 2385 1650
rect 3210 1710 3590 1720
rect 3210 1630 3220 1710
rect 3580 1630 3590 1710
rect 3210 1620 3590 1630
rect -790 1585 -10 1595
rect -790 25 -780 1585
rect -420 25 -380 1585
rect -20 25 -10 1585
rect -790 15 -10 25
rect -390 -20 -10 15
rect -390 -100 -380 -20
rect -20 -100 -10 -20
rect -390 -110 -10 -100
rect 410 1585 790 1595
rect 410 25 420 1585
rect 780 25 790 1585
rect 410 -20 790 25
rect 1210 1585 1590 1595
rect 1210 25 1220 1585
rect 1580 25 1590 1585
rect 1210 15 1590 25
rect 2010 1585 2390 1595
rect 2010 25 2020 1585
rect 2380 25 2390 1585
rect 410 -100 420 -20
rect 780 -100 790 -20
rect 410 -110 790 -100
rect 1215 -380 1585 -370
rect 1215 -455 1225 -380
rect 1575 -455 1585 -380
rect 1215 -465 1585 -455
rect -790 -815 -10 -805
rect -790 -2375 -780 -815
rect -420 -2375 -380 -815
rect -20 -2375 -10 -815
rect -790 -2385 -10 -2375
rect -390 -2420 -10 -2385
rect -390 -2500 -380 -2420
rect -20 -2500 -10 -2420
rect -390 -2510 -10 -2500
rect 410 -815 790 -805
rect 410 -2375 420 -815
rect 780 -2375 790 -815
rect 410 -2420 790 -2375
rect 1210 -815 1590 -805
rect 1210 -2375 1220 -815
rect 1580 -2375 1590 -815
rect 1210 -2385 1590 -2375
rect 2010 -815 2390 25
rect 2010 -2375 2020 -815
rect 2380 -2375 2390 -815
rect 2010 -2385 2390 -2375
rect 2810 1585 3190 1595
rect 2810 25 2820 1585
rect 3180 25 3190 1585
rect 2810 -815 3190 25
rect 3610 1585 3990 1795
rect 5215 1725 5585 1735
rect 5215 1650 5225 1725
rect 5575 1650 5585 1725
rect 8415 1725 8785 1735
rect 5215 1640 5585 1650
rect 7210 1710 7590 1720
rect 7210 1630 7220 1710
rect 7580 1630 7590 1710
rect 8415 1650 8425 1725
rect 8775 1650 8785 1725
rect 8415 1640 8785 1650
rect 14015 1725 14385 1735
rect 14015 1650 14025 1725
rect 14375 1650 14385 1725
rect 14015 1640 14385 1650
rect 20015 1725 20385 1735
rect 20015 1650 20025 1725
rect 20375 1650 20385 1725
rect 20015 1640 20385 1650
rect 21615 1725 21985 1735
rect 21615 1650 21625 1725
rect 21975 1650 21985 1725
rect 21615 1640 21985 1650
rect 7210 1620 7590 1630
rect 3610 25 3620 1585
rect 3980 25 3990 1585
rect 3610 15 3990 25
rect 4410 1585 4790 1595
rect 4410 25 4420 1585
rect 4780 25 4790 1585
rect 3630 -365 4000 -355
rect 3630 -440 3640 -365
rect 3990 -440 4000 -365
rect 3630 -450 4000 -440
rect 3210 -690 3590 -680
rect 3210 -770 3220 -690
rect 3580 -770 3590 -690
rect 3210 -780 3590 -770
rect 2810 -2375 2820 -815
rect 3180 -2375 3190 -815
rect 410 -2500 420 -2420
rect 780 -2500 790 -2420
rect 410 -2510 790 -2500
rect 2015 -2440 2385 -2430
rect 2015 -2515 2025 -2440
rect 2375 -2515 2385 -2440
rect 2015 -2525 2385 -2515
rect 2015 -3195 2385 -3185
rect 2015 -3270 2025 -3195
rect 2375 -3270 2385 -3195
rect 2015 -3280 2385 -3270
rect -790 -3335 -10 -3325
rect -790 -4895 -780 -3335
rect -420 -4895 -380 -3335
rect -20 -4895 -10 -3335
rect -790 -4905 -10 -4895
rect -390 -4940 -10 -4905
rect -390 -5020 -380 -4940
rect -20 -5020 -10 -4940
rect -390 -5030 -10 -5020
rect 410 -3335 790 -3325
rect 410 -4895 420 -3335
rect 780 -4895 790 -3335
rect 410 -5270 790 -4895
rect 1210 -3335 1590 -3325
rect 1210 -4895 1220 -3335
rect 1580 -4895 1590 -3335
rect 1210 -5005 1590 -4895
rect 1210 -5085 1220 -5005
rect 1580 -5085 1590 -5005
rect 1210 -5095 1590 -5085
rect 2010 -3335 2390 -3325
rect 2010 -4895 2020 -3335
rect 2380 -4895 2390 -3335
rect 1215 -5145 1585 -5135
rect 1215 -5220 1225 -5145
rect 1575 -5220 1585 -5145
rect 1215 -5230 1585 -5220
rect 2010 -5270 2390 -4895
rect 2810 -3335 3190 -2375
rect 3610 -815 3990 -805
rect 3610 -2375 3620 -815
rect 3980 -2375 3990 -815
rect 3610 -2460 3990 -2375
rect 4410 -815 4790 25
rect 5210 1585 5590 1595
rect 5210 25 5220 1585
rect 5580 25 5590 1585
rect 5210 15 5590 25
rect 6010 1585 6390 1595
rect 6010 25 6020 1585
rect 6380 25 6390 1585
rect 5820 -20 5990 -10
rect 5820 -80 5830 -20
rect 5980 -80 5990 -20
rect 5820 -90 5990 -80
rect 5220 -380 5590 -370
rect 5220 -455 5230 -380
rect 5580 -455 5590 -380
rect 5220 -465 5590 -455
rect 5820 -710 5990 -700
rect 5820 -770 5830 -710
rect 5980 -770 5990 -710
rect 5820 -780 5990 -770
rect 4410 -2375 4420 -815
rect 4780 -2375 4790 -815
rect 4410 -2385 4790 -2375
rect 5210 -815 5590 -805
rect 5210 -2375 5220 -815
rect 5580 -2375 5590 -815
rect 5210 -2385 5590 -2375
rect 6010 -815 6390 25
rect 6810 1585 7190 1595
rect 6810 25 6820 1585
rect 7180 25 7190 1585
rect 6410 -20 6580 -10
rect 6410 -80 6420 -20
rect 6570 -80 6580 -20
rect 6410 -90 6580 -80
rect 6810 -125 7190 25
rect 6810 -205 6820 -125
rect 7180 -205 7190 -125
rect 6410 -710 6580 -700
rect 6410 -770 6420 -710
rect 6570 -770 6580 -710
rect 6410 -780 6580 -770
rect 6010 -2375 6020 -815
rect 6380 -2375 6390 -815
rect 6010 -2385 6390 -2375
rect 6810 -815 7190 -205
rect 7610 1585 7990 1595
rect 7610 25 7620 1585
rect 7980 25 7990 1585
rect 7210 -690 7590 -680
rect 7210 -770 7220 -690
rect 7580 -770 7590 -690
rect 7210 -780 7590 -770
rect 6810 -2375 6820 -815
rect 7180 -2375 7190 -815
rect 3610 -2540 3620 -2460
rect 3980 -2540 3990 -2460
rect 5215 -2440 5585 -2430
rect 5215 -2515 5225 -2440
rect 5575 -2515 5585 -2440
rect 5215 -2525 5585 -2515
rect 3610 -2550 3990 -2540
rect 6810 -2710 7190 -2375
rect 6810 -2790 6820 -2710
rect 7180 -2790 7190 -2710
rect 4410 -3190 4790 -3180
rect 6010 -3185 6390 -3175
rect 4410 -3270 4420 -3190
rect 4780 -3270 4790 -3190
rect 2810 -4895 2820 -3335
rect 3180 -4895 3190 -3335
rect 2810 -5005 3190 -4895
rect 2810 -5085 2820 -5005
rect 3180 -5085 3190 -5005
rect 2810 -5095 3190 -5085
rect 3610 -3335 3990 -3325
rect 3610 -4895 3620 -3335
rect 3980 -4895 3990 -3335
rect 3610 -5270 3990 -4895
rect 4410 -3335 4790 -3270
rect 5215 -3195 5585 -3185
rect 5215 -3270 5225 -3195
rect 5575 -3270 5585 -3195
rect 5215 -3280 5585 -3270
rect 6010 -3265 6020 -3185
rect 6380 -3265 6390 -3185
rect 4410 -4895 4420 -3335
rect 4780 -4895 4790 -3335
rect 4410 -4930 4790 -4895
rect 5210 -3335 5590 -3325
rect 5210 -4895 5220 -3335
rect 5580 -4895 5590 -3335
rect 4410 -4940 4450 -4930
rect 4410 -4960 4420 -4940
rect 4440 -4960 4450 -4940
rect 4410 -4970 4450 -4960
rect -795 -5370 3990 -5270
rect -790 -5735 -10 -5725
rect -790 -7295 -780 -5735
rect -420 -7295 -380 -5735
rect -20 -7295 -10 -5735
rect -790 -7305 -10 -7295
rect 410 -5735 790 -5370
rect 410 -7295 420 -5735
rect 780 -7295 790 -5735
rect 410 -7305 790 -7295
rect 1210 -5545 1590 -5535
rect 1210 -5625 1220 -5545
rect 1580 -5625 1590 -5545
rect 1210 -5735 1590 -5625
rect 1210 -7295 1220 -5735
rect 1580 -7295 1590 -5735
rect 1210 -7305 1590 -7295
rect 2010 -5735 2390 -5370
rect 2010 -7295 2020 -5735
rect 2380 -7295 2390 -5735
rect 2010 -7305 2390 -7295
rect 2810 -5545 3190 -5535
rect 2810 -5625 2820 -5545
rect 3180 -5625 3190 -5545
rect 2810 -5735 3190 -5625
rect 2810 -7295 2820 -5735
rect 3180 -7295 3190 -5735
rect 2810 -7305 3190 -7295
rect 3610 -5735 3990 -5370
rect 4415 -5140 4785 -5130
rect 4415 -5490 4425 -5140
rect 4775 -5490 4785 -5140
rect 4415 -5500 4785 -5490
rect 3610 -7295 3620 -5735
rect 3980 -7295 3990 -5735
rect 3610 -7305 3990 -7295
rect 4410 -5670 4450 -5660
rect 4410 -5690 4420 -5670
rect 4440 -5690 4450 -5670
rect 4410 -5700 4450 -5690
rect 4410 -5735 4790 -5700
rect 4410 -7295 4420 -5735
rect 4780 -7295 4790 -5735
rect -390 -7340 -10 -7305
rect -390 -7420 -380 -7340
rect -20 -7420 -10 -7340
rect -390 -7430 -10 -7420
rect 2015 -7360 2385 -7350
rect 2015 -7435 2025 -7360
rect 2375 -7435 2385 -7360
rect 2015 -7445 2385 -7435
rect 3615 -7360 3985 -7350
rect 3615 -7435 3625 -7360
rect 3975 -7435 3985 -7360
rect 3615 -7445 3985 -7435
rect 4410 -7360 4790 -7295
rect 5210 -5735 5590 -4895
rect 5210 -7295 5220 -5735
rect 5580 -7295 5590 -5735
rect 5210 -7305 5590 -7295
rect 6010 -3335 6390 -3265
rect 6010 -4895 6020 -3335
rect 6380 -4895 6390 -3335
rect 6010 -5735 6390 -4895
rect 6810 -3335 7190 -2790
rect 7610 -815 7990 25
rect 8410 1585 8790 1595
rect 8410 25 8420 1585
rect 8780 25 8790 1585
rect 8020 -440 8390 -430
rect 8020 -515 8030 -440
rect 8380 -515 8390 -440
rect 8020 -525 8390 -515
rect 7610 -2375 7620 -815
rect 7980 -2375 7990 -815
rect 7610 -3260 7990 -2375
rect 8410 -815 8790 25
rect 9210 1585 9590 1595
rect 9210 25 9220 1585
rect 9580 25 9590 1585
rect 9210 15 9590 25
rect 10010 1585 10390 1595
rect 10010 25 10020 1585
rect 10380 25 10390 1585
rect 10010 -20 10390 25
rect 10010 -100 10020 -20
rect 10380 -100 10390 -20
rect 10010 -110 10390 -100
rect 10810 1585 11990 1595
rect 10810 25 10820 1585
rect 11180 25 11220 1585
rect 11580 25 11620 1585
rect 11980 25 11990 1585
rect 10810 15 11990 25
rect 10810 -20 11190 15
rect 10810 -100 10820 -20
rect 11180 -100 11190 -20
rect 10810 -110 11190 -100
rect 11610 -20 11990 15
rect 11610 -100 11620 -20
rect 11980 -100 11990 -20
rect 11610 -110 11990 -100
rect 12410 1585 12790 1595
rect 12410 25 12420 1585
rect 12780 25 12790 1585
rect 12410 -665 12790 25
rect 12410 -745 12420 -665
rect 12780 -745 12790 -665
rect 8410 -2375 8420 -815
rect 8780 -2375 8790 -815
rect 8410 -2385 8790 -2375
rect 9210 -815 9590 -805
rect 9210 -2375 9220 -815
rect 9580 -2375 9590 -815
rect 9210 -2385 9590 -2375
rect 10010 -815 10390 -805
rect 10010 -2375 10020 -815
rect 10380 -2375 10390 -815
rect 10010 -2420 10390 -2375
rect 8415 -2440 8785 -2430
rect 8415 -2515 8425 -2440
rect 8775 -2515 8785 -2440
rect 10010 -2500 10020 -2420
rect 10380 -2500 10390 -2420
rect 10010 -2510 10390 -2500
rect 10810 -815 11990 -805
rect 10810 -2375 10820 -815
rect 11180 -2375 11220 -815
rect 11580 -2375 11620 -815
rect 11980 -2375 11990 -815
rect 10810 -2385 11990 -2375
rect 10810 -2420 11190 -2385
rect 10810 -2500 10820 -2420
rect 11180 -2500 11190 -2420
rect 10810 -2510 11190 -2500
rect 11610 -2420 11990 -2385
rect 11610 -2500 11620 -2420
rect 11980 -2500 11990 -2420
rect 11610 -2510 11990 -2500
rect 12410 -815 12790 -745
rect 12410 -2375 12420 -815
rect 12780 -2375 12790 -815
rect 8415 -2525 8785 -2515
rect 7560 -3270 7990 -3260
rect 7560 -3290 7570 -3270
rect 7590 -3290 7990 -3270
rect 8415 -3195 8785 -3185
rect 8415 -3270 8425 -3195
rect 8775 -3270 8785 -3195
rect 8415 -3280 8785 -3270
rect 7560 -3300 7990 -3290
rect 6810 -4895 6820 -3335
rect 7180 -4895 7190 -3335
rect 6410 -4940 6790 -4930
rect 6410 -5025 6420 -4940
rect 6780 -5025 6790 -4940
rect 6410 -5035 6790 -5025
rect 6415 -5140 6785 -5130
rect 6415 -5490 6425 -5140
rect 6775 -5490 6785 -5140
rect 6415 -5500 6785 -5490
rect 6410 -5605 6790 -5595
rect 6410 -5690 6420 -5605
rect 6780 -5690 6790 -5605
rect 6410 -5700 6790 -5690
rect 6010 -7295 6020 -5735
rect 6380 -7295 6390 -5735
rect 6010 -7305 6390 -7295
rect 6810 -5735 7190 -4895
rect 6810 -7295 6820 -5735
rect 7180 -7295 7190 -5735
rect 6810 -7305 7190 -7295
rect 7610 -3335 7990 -3325
rect 7610 -4895 7620 -3335
rect 7980 -4895 7990 -3335
rect 7610 -5735 7990 -4895
rect 8410 -3335 8790 -3325
rect 8410 -4895 8420 -3335
rect 8780 -4895 8790 -3335
rect 8410 -4905 8790 -4895
rect 9210 -3335 9590 -3325
rect 9210 -4895 9220 -3335
rect 9580 -4895 9590 -3335
rect 8415 -5140 8785 -5130
rect 8415 -5490 8425 -5140
rect 8775 -5490 8785 -5140
rect 8415 -5500 8785 -5490
rect 7610 -7295 7620 -5735
rect 7980 -7295 7990 -5735
rect 7610 -7305 7990 -7295
rect 8410 -5735 8790 -5725
rect 8410 -7295 8420 -5735
rect 8780 -7295 8790 -5735
rect 8410 -7305 8790 -7295
rect 9210 -5735 9590 -4895
rect 9210 -7295 9220 -5735
rect 9580 -7295 9590 -5735
rect 9210 -7305 9590 -7295
rect 10010 -3335 10390 -3325
rect 10010 -4895 10020 -3335
rect 10380 -4895 10390 -3335
rect 10010 -5645 10390 -4895
rect 10810 -3335 11990 -3325
rect 10810 -4895 10820 -3335
rect 11180 -4895 11220 -3335
rect 11580 -4895 11620 -3335
rect 11980 -4895 11990 -3335
rect 10810 -4905 11990 -4895
rect 10810 -4940 11190 -4905
rect 10810 -5020 10820 -4940
rect 11180 -5020 11190 -4940
rect 10810 -5030 11190 -5020
rect 11610 -4940 11990 -4905
rect 11610 -5020 11620 -4940
rect 11980 -5020 11990 -4940
rect 11610 -5030 11990 -5020
rect 12410 -3335 12790 -2375
rect 13210 1585 13590 1595
rect 13210 25 13220 1585
rect 13580 25 13590 1585
rect 13210 -815 13590 25
rect 14010 1585 14390 1595
rect 14010 25 14020 1585
rect 14380 25 14390 1585
rect 14010 10 14390 25
rect 14810 1585 15190 1595
rect 14810 25 14820 1585
rect 15180 25 15190 1585
rect 14015 -250 14385 -240
rect 14015 -325 14025 -250
rect 14375 -325 14385 -250
rect 14015 -335 14385 -325
rect 13210 -2375 13220 -815
rect 13580 -2375 13590 -815
rect 13210 -2385 13590 -2375
rect 14010 -815 14390 -800
rect 14010 -2375 14020 -815
rect 14380 -2375 14390 -815
rect 14010 -2385 14390 -2375
rect 14810 -815 15190 25
rect 14810 -2375 14820 -815
rect 15180 -2375 15190 -815
rect 14810 -2385 15190 -2375
rect 15610 1585 15990 1595
rect 15610 25 15620 1585
rect 15980 25 15990 1585
rect 15610 -815 15990 25
rect 16410 1585 17190 1595
rect 16410 25 16420 1585
rect 16780 25 16820 1585
rect 17180 25 17190 1585
rect 16410 15 17190 25
rect 18010 1585 18790 1595
rect 18010 25 18020 1585
rect 18380 25 18420 1585
rect 18780 25 18790 1585
rect 18010 15 18790 25
rect 19210 1585 19590 1595
rect 19210 25 19220 1585
rect 19580 25 19590 1585
rect 19210 15 19590 25
rect 20010 1585 20390 1595
rect 20010 25 20020 1585
rect 20380 25 20390 1585
rect 20010 15 20390 25
rect 20810 1585 21190 1595
rect 20810 25 20820 1585
rect 21180 25 21190 1585
rect 20810 15 21190 25
rect 21610 1585 21990 1595
rect 21610 25 21620 1585
rect 21980 25 21990 1585
rect 21610 15 21990 25
rect 22410 1585 22790 1595
rect 22410 25 22420 1585
rect 22780 25 22790 1585
rect 22410 15 22790 25
rect 23210 1585 23990 1595
rect 23210 25 23220 1585
rect 23580 25 23620 1585
rect 23980 25 23990 1585
rect 23210 15 23990 25
rect 16410 -20 16790 15
rect 16410 -100 16420 -20
rect 16780 -100 16790 -20
rect 16410 -110 16790 -100
rect 18410 -20 18790 15
rect 18410 -100 18420 -20
rect 18780 -100 18790 -20
rect 18410 -110 18790 -100
rect 20200 -35 20390 15
rect 21610 -35 21800 15
rect 20200 -135 21800 -35
rect 23210 -20 23590 15
rect 23210 -100 23220 -20
rect 23580 -100 23590 -20
rect 23210 -110 23590 -100
rect 21625 -385 21995 -375
rect 20015 -400 20385 -390
rect 20015 -475 20025 -400
rect 20375 -475 20385 -400
rect 21625 -460 21635 -385
rect 21985 -460 21995 -385
rect 21625 -470 21995 -460
rect 20015 -485 20385 -475
rect 20200 -755 21800 -655
rect 20200 -805 20390 -755
rect 21610 -805 21800 -755
rect 15610 -2375 15620 -815
rect 15980 -2375 15990 -815
rect 14015 -2440 14385 -2430
rect 14015 -2515 14025 -2440
rect 14375 -2515 14385 -2440
rect 14015 -2525 14385 -2515
rect 15610 -2960 15990 -2375
rect 16410 -815 17190 -805
rect 16410 -2375 16420 -815
rect 16780 -2375 16820 -815
rect 17180 -2375 17190 -815
rect 16410 -2385 17190 -2375
rect 18010 -815 18790 -805
rect 18010 -2375 18020 -815
rect 18380 -2375 18420 -815
rect 18780 -2375 18790 -815
rect 18010 -2385 18790 -2375
rect 19210 -815 19590 -805
rect 19210 -2375 19220 -815
rect 19580 -2375 19590 -815
rect 19210 -2385 19590 -2375
rect 20010 -815 20390 -805
rect 20010 -2375 20020 -815
rect 20380 -2375 20390 -815
rect 20010 -2385 20390 -2375
rect 20810 -815 21190 -805
rect 20810 -2375 20820 -815
rect 21180 -2375 21190 -815
rect 20810 -2385 21190 -2375
rect 21610 -815 21990 -805
rect 21610 -2375 21620 -815
rect 21980 -2375 21990 -815
rect 21610 -2385 21990 -2375
rect 22410 -815 22790 -805
rect 22410 -2375 22420 -815
rect 22780 -2375 22790 -815
rect 22410 -2385 22790 -2375
rect 23210 -815 23990 -805
rect 23210 -2375 23220 -815
rect 23580 -2375 23620 -815
rect 23980 -2375 23990 -815
rect 23210 -2385 23990 -2375
rect 16410 -2420 16790 -2385
rect 16410 -2500 16420 -2420
rect 16780 -2500 16790 -2420
rect 16410 -2510 16790 -2500
rect 18410 -2420 18790 -2385
rect 18410 -2500 18420 -2420
rect 18780 -2500 18790 -2420
rect 18410 -2510 18790 -2500
rect 23210 -2420 23590 -2385
rect 23210 -2500 23220 -2420
rect 23580 -2500 23590 -2420
rect 23210 -2510 23590 -2500
rect 21615 -2765 21985 -2755
rect 20015 -2780 20385 -2770
rect 20015 -2855 20025 -2780
rect 20375 -2855 20385 -2780
rect 21615 -2840 21625 -2765
rect 21975 -2840 21985 -2765
rect 21615 -2850 21985 -2840
rect 20015 -2865 20385 -2855
rect 15610 -2970 23950 -2960
rect 15610 -3050 19610 -2970
rect 19990 -3050 20410 -2970
rect 20790 -3050 21210 -2970
rect 21590 -3050 22010 -2970
rect 22390 -3050 23950 -2970
rect 15610 -3060 23950 -3050
rect 14015 -3190 14385 -3180
rect 14015 -3265 14025 -3190
rect 14375 -3265 14385 -3190
rect 14015 -3275 14385 -3265
rect 12410 -4895 12420 -3335
rect 12780 -4895 12790 -3335
rect 10010 -5665 10020 -5645
rect 10040 -5665 10390 -5645
rect 10010 -5735 10390 -5665
rect 10010 -7295 10020 -5735
rect 10380 -7295 10390 -5735
rect 10010 -7305 10390 -7295
rect 10810 -5735 11990 -5725
rect 10810 -7295 10820 -5735
rect 11180 -7295 11220 -5735
rect 11580 -7295 11620 -5735
rect 11980 -7295 11990 -5735
rect 10810 -7305 11990 -7295
rect 12410 -5735 12790 -4895
rect 12410 -7295 12420 -5735
rect 12780 -7295 12790 -5735
rect 12410 -7305 12790 -7295
rect 13210 -3335 13590 -3325
rect 13210 -4895 13220 -3335
rect 13580 -4895 13590 -3335
rect 13210 -5735 13590 -4895
rect 14010 -3335 14390 -3325
rect 14010 -4895 14020 -3335
rect 14380 -4895 14390 -3335
rect 14010 -4910 14390 -4895
rect 14810 -3335 15190 -3325
rect 14810 -4895 14820 -3335
rect 15180 -4895 15190 -3335
rect 14015 -5180 14385 -5170
rect 14015 -5530 14025 -5180
rect 14375 -5530 14385 -5180
rect 14015 -5540 14385 -5530
rect 13210 -7295 13220 -5735
rect 13580 -7295 13590 -5735
rect 13210 -7305 13590 -7295
rect 14010 -5735 14390 -5720
rect 14010 -7295 14015 -5735
rect 14380 -7295 14390 -5735
rect 14010 -7305 14390 -7295
rect 14810 -5735 15190 -4895
rect 14810 -7295 14820 -5735
rect 15180 -7295 15190 -5735
rect 14810 -7305 15190 -7295
rect 15610 -3335 15990 -3060
rect 20200 -3275 21800 -3175
rect 20200 -3325 20390 -3275
rect 21610 -3325 21800 -3275
rect 15610 -4895 15620 -3335
rect 15980 -4895 15990 -3335
rect 15610 -5735 15990 -4895
rect 16410 -3335 17190 -3325
rect 16410 -4895 16420 -3335
rect 16780 -4895 16820 -3335
rect 17180 -4895 17190 -3335
rect 16410 -4905 17190 -4895
rect 18010 -3335 18790 -3325
rect 18010 -4895 18020 -3335
rect 18380 -4895 18420 -3335
rect 18780 -4895 18790 -3335
rect 18010 -4905 18790 -4895
rect 19210 -3335 19590 -3325
rect 19210 -4895 19220 -3335
rect 19580 -4895 19590 -3335
rect 19210 -4905 19590 -4895
rect 20010 -3335 20390 -3325
rect 20010 -4895 20020 -3335
rect 20380 -4895 20390 -3335
rect 20010 -4905 20390 -4895
rect 20810 -3335 21190 -3325
rect 20810 -4895 20820 -3335
rect 21180 -4895 21190 -3335
rect 20810 -4905 21190 -4895
rect 21610 -3335 21990 -3325
rect 21610 -4895 21620 -3335
rect 21980 -4895 21990 -3335
rect 21610 -4905 21990 -4895
rect 22410 -3335 22790 -3325
rect 22410 -4895 22420 -3335
rect 22780 -4895 22790 -3335
rect 22410 -4905 22790 -4895
rect 23210 -3335 23990 -3325
rect 23210 -4895 23220 -3335
rect 23580 -4895 23620 -3335
rect 23980 -4895 23990 -3335
rect 23210 -4905 23990 -4895
rect 16410 -4940 16790 -4905
rect 16410 -5020 16420 -4940
rect 16780 -5020 16790 -4940
rect 16410 -5030 16790 -5020
rect 18410 -4940 18790 -4905
rect 18410 -5020 18420 -4940
rect 18780 -5020 18790 -4940
rect 18410 -5030 18790 -5020
rect 23210 -4940 23590 -4905
rect 23210 -5020 23220 -4940
rect 23580 -5020 23590 -4940
rect 23210 -5030 23590 -5020
rect 19270 -5095 19640 -5085
rect 19270 -5445 19280 -5095
rect 19630 -5445 19640 -5095
rect 22330 -5110 22700 -5100
rect 19270 -5455 19640 -5445
rect 20200 -5520 21800 -5420
rect 22330 -5460 22340 -5110
rect 22690 -5460 22700 -5110
rect 22330 -5470 22700 -5460
rect 20200 -5725 20390 -5520
rect 15610 -7295 15620 -5735
rect 15980 -7295 15990 -5735
rect 15610 -7305 15990 -7295
rect 16410 -5735 17190 -5725
rect 16410 -7295 16420 -5735
rect 16780 -7295 16820 -5735
rect 17180 -7295 17190 -5735
rect 16410 -7305 17190 -7295
rect 18010 -5735 18790 -5725
rect 18010 -7295 18020 -5735
rect 18380 -7295 18420 -5735
rect 18010 -7300 18420 -7295
rect 18780 -7300 18790 -5735
rect 18010 -7305 18790 -7300
rect 19210 -5735 19590 -5725
rect 19210 -7295 19220 -5735
rect 19580 -7295 19590 -5735
rect 19210 -7305 19590 -7295
rect 20010 -5735 20390 -5725
rect 20010 -7295 20020 -5735
rect 20380 -7295 20390 -5735
rect 20010 -7305 20390 -7295
rect 20810 -5555 21190 -5545
rect 20810 -5635 20820 -5555
rect 21180 -5635 21190 -5555
rect 20810 -5735 21190 -5635
rect 20810 -7295 20820 -5735
rect 21180 -7295 21190 -5735
rect 20810 -7305 21190 -7295
rect 21610 -5725 21800 -5520
rect 21610 -5735 21990 -5725
rect 21610 -7295 21620 -5735
rect 21980 -7295 21990 -5735
rect 21610 -7305 21990 -7295
rect 22410 -5735 22790 -5725
rect 22410 -7295 22420 -5735
rect 22780 -7295 22790 -5735
rect 22410 -7305 22790 -7295
rect 23210 -5735 23990 -5725
rect 23210 -7295 23220 -5735
rect 23580 -7295 23620 -5735
rect 23980 -7295 23990 -5735
rect 23210 -7305 23990 -7295
rect 7200 -7340 7600 -7330
rect 4410 -7440 4420 -7360
rect 4780 -7440 4790 -7360
rect 4410 -7450 4790 -7440
rect 6015 -7360 6385 -7350
rect 6015 -7435 6025 -7360
rect 6375 -7435 6385 -7360
rect 6015 -7445 6385 -7435
rect 7200 -7420 7210 -7340
rect 7590 -7420 7600 -7340
rect 7200 -7455 7600 -7420
rect 8000 -7340 8400 -7330
rect 8000 -7420 8010 -7340
rect 8390 -7420 8400 -7340
rect 8000 -7455 8400 -7420
rect 8420 -7360 8780 -7305
rect 8420 -7425 8430 -7360
rect 8770 -7425 8780 -7360
rect 8420 -7435 8780 -7425
rect 8800 -7340 9200 -7330
rect 8800 -7420 8810 -7340
rect 9190 -7420 9200 -7340
rect 8800 -7455 9200 -7420
rect 9600 -7340 10000 -7330
rect 9600 -7420 9610 -7340
rect 9990 -7420 10000 -7340
rect 9600 -7455 10000 -7420
rect 10810 -7340 11190 -7305
rect 10810 -7420 10820 -7340
rect 11180 -7420 11190 -7340
rect 10810 -7430 11190 -7420
rect 11610 -7340 11990 -7305
rect 11610 -7420 11620 -7340
rect 11980 -7420 11990 -7340
rect 11610 -7430 11990 -7420
rect 12800 -7340 13200 -7330
rect 12800 -7420 12810 -7340
rect 13190 -7420 13200 -7340
rect 12800 -7455 13200 -7420
rect 13600 -7340 14000 -7330
rect 13600 -7420 13610 -7340
rect 13990 -7420 14000 -7340
rect 13600 -7455 14000 -7420
rect 14020 -7360 14380 -7305
rect 14020 -7425 14030 -7360
rect 14370 -7425 14380 -7360
rect 14020 -7435 14380 -7425
rect 16410 -7340 16790 -7305
rect 16410 -7420 16420 -7340
rect 16780 -7420 16790 -7340
rect 16410 -7430 16790 -7420
rect 18410 -7340 18790 -7305
rect 18410 -7420 18420 -7340
rect 18780 -7420 18790 -7340
rect 18410 -7430 18790 -7420
rect 19600 -7340 20000 -7330
rect 19600 -7420 19610 -7340
rect 19990 -7420 20000 -7340
rect 19600 -7455 20000 -7420
rect 20400 -7340 20800 -7330
rect 20400 -7420 20410 -7340
rect 20790 -7420 20800 -7340
rect 21200 -7340 21600 -7330
rect 20400 -7455 20800 -7420
rect 20820 -7360 21180 -7350
rect 20820 -7425 20830 -7360
rect 21170 -7425 21180 -7360
rect 20820 -7435 21180 -7425
rect 21200 -7420 21210 -7340
rect 21590 -7420 21600 -7340
rect 21200 -7455 21600 -7420
rect 22000 -7340 22400 -7330
rect 22000 -7420 22010 -7340
rect 22390 -7420 22400 -7340
rect 22000 -7455 22400 -7420
rect 23210 -7340 23590 -7305
rect 23210 -7420 23220 -7340
rect 23580 -7420 23590 -7340
rect 23210 -7430 23590 -7420
rect 7200 -7555 24030 -7455
<< viali >>
rect 2025 1650 2375 1725
rect 3220 1630 3580 1710
rect -780 25 -420 1585
rect -380 25 -20 1585
rect 1220 25 1580 1585
rect 1225 -455 1575 -380
rect -780 -2375 -420 -815
rect -380 -2375 -20 -815
rect 1220 -2375 1580 -815
rect 5225 1650 5575 1725
rect 7220 1630 7580 1710
rect 8425 1650 8775 1725
rect 14025 1650 14375 1725
rect 20025 1650 20375 1725
rect 21625 1650 21975 1725
rect 3640 -440 3990 -365
rect 3220 -770 3580 -690
rect 2025 -2515 2375 -2440
rect 2025 -3270 2375 -3195
rect -780 -4895 -420 -3335
rect -380 -4895 -20 -3335
rect 1225 -5220 1575 -5145
rect 5220 25 5580 1585
rect 5830 -80 5980 -20
rect 5230 -455 5580 -380
rect 5830 -770 5980 -710
rect 5220 -2375 5580 -815
rect 6420 -80 6570 -20
rect 6420 -770 6570 -710
rect 7220 -770 7580 -690
rect 5225 -2515 5575 -2440
rect 5225 -3270 5575 -3195
rect 6020 -3265 6380 -3185
rect 4420 -4895 4780 -3335
rect -780 -7295 -420 -5735
rect -380 -7295 -20 -5735
rect 4425 -5490 4775 -5140
rect 4420 -7295 4780 -5735
rect 2025 -7435 2375 -7360
rect 3625 -7435 3975 -7360
rect 8030 -515 8380 -440
rect 9220 25 9580 1585
rect 10020 25 10380 1585
rect 10820 25 11180 1585
rect 11220 25 11580 1585
rect 11620 25 11980 1585
rect 9220 -2375 9580 -815
rect 10020 -2375 10380 -815
rect 8425 -2515 8775 -2440
rect 10820 -2375 11180 -815
rect 11220 -2375 11580 -815
rect 11620 -2375 11980 -815
rect 8425 -3270 8775 -3195
rect 6420 -5025 6780 -4940
rect 6425 -5490 6775 -5140
rect 6420 -5690 6780 -5605
rect 8420 -4895 8780 -3335
rect 8425 -5490 8775 -5140
rect 8420 -7295 8780 -5735
rect 10820 -4895 11180 -3335
rect 11220 -4895 11580 -3335
rect 11620 -4895 11980 -3335
rect 14020 25 14380 1585
rect 14025 -325 14375 -250
rect 14020 -2375 14380 -815
rect 16420 25 16780 1585
rect 16820 25 17180 1585
rect 18020 25 18380 1585
rect 18420 25 18780 1585
rect 19220 25 19580 1585
rect 20820 25 21180 1585
rect 22420 25 22780 1585
rect 23220 25 23580 1585
rect 23620 25 23980 1585
rect 20025 -475 20375 -400
rect 21635 -460 21985 -385
rect 14025 -2515 14375 -2440
rect 16420 -2375 16780 -815
rect 16820 -2375 17180 -815
rect 18020 -2375 18380 -815
rect 18420 -2375 18780 -815
rect 19220 -2375 19580 -815
rect 20820 -2375 21180 -815
rect 22420 -2375 22780 -815
rect 23220 -2375 23580 -815
rect 23620 -2375 23980 -815
rect 20025 -2855 20375 -2780
rect 21625 -2840 21975 -2765
rect 14025 -3265 14375 -3190
rect 10820 -7295 11180 -5735
rect 11220 -7295 11580 -5735
rect 11620 -7295 11980 -5735
rect 14020 -4895 14380 -3335
rect 14025 -5530 14375 -5180
rect 14015 -7295 14380 -5735
rect 16420 -4895 16780 -3335
rect 16820 -4895 17180 -3335
rect 18020 -4895 18380 -3335
rect 18420 -4895 18780 -3335
rect 19220 -4895 19580 -3335
rect 20820 -4895 21180 -3335
rect 22420 -4895 22780 -3335
rect 23220 -4895 23580 -3335
rect 23620 -4895 23980 -3335
rect 19280 -5445 19630 -5095
rect 22340 -5460 22690 -5110
rect 16420 -7295 16780 -5735
rect 16820 -7295 17180 -5735
rect 18020 -7295 18380 -5735
rect 18420 -7300 18780 -5740
rect 19220 -7295 19580 -5735
rect 20820 -7295 21180 -5735
rect 22420 -7295 22780 -5735
rect 23220 -7295 23580 -5735
rect 23620 -7295 23980 -5735
rect 6025 -7435 6375 -7360
rect 8430 -7425 8770 -7360
rect 20830 -7425 21170 -7360
<< metal1 >>
rect 20075 2595 21945 2600
rect -800 1900 24000 2595
rect -800 1725 19600 1900
rect -800 1650 2025 1725
rect 2375 1710 5225 1725
rect 2375 1650 3220 1710
rect -800 1630 3220 1650
rect 3580 1650 5225 1710
rect 5575 1710 8425 1725
rect 5575 1650 7220 1710
rect 3580 1630 7220 1650
rect 7580 1650 8425 1710
rect 8775 1650 14025 1725
rect 14375 1650 19600 1725
rect 7580 1635 19600 1650
rect 7580 1630 17590 1635
rect -800 1595 17590 1630
rect -800 1585 5785 1595
rect -800 25 -780 1585
rect -420 25 -380 1585
rect -20 25 1220 1585
rect 1580 25 5220 1585
rect 5580 25 5785 1585
rect -800 -365 5785 25
rect 6610 1585 17590 1595
rect 6610 25 9220 1585
rect 9580 25 10020 1585
rect 10380 25 10820 1585
rect 11180 25 11220 1585
rect 11580 25 11620 1585
rect 11980 25 14020 1585
rect 14380 25 16420 1585
rect 16780 25 16820 1585
rect 17180 25 17590 1585
rect 5930 -10 6470 5
rect 5820 -20 6580 -10
rect 5820 -80 5830 -20
rect 5980 -80 6420 -20
rect 6570 -80 6580 -20
rect 5820 -90 6580 -80
rect -800 -380 3640 -365
rect -800 -455 1225 -380
rect 1575 -440 3640 -380
rect 3990 -380 5785 -365
rect 3990 -440 5230 -380
rect 1575 -455 5230 -440
rect 5580 -455 5785 -380
rect -800 -690 5785 -455
rect -800 -770 3220 -690
rect 3580 -770 5785 -690
rect 5930 -700 6470 -90
rect 6610 -250 17590 25
rect 6610 -325 14025 -250
rect 14375 -325 17590 -250
rect 6610 -440 17590 -325
rect 6610 -515 8030 -440
rect 8380 -515 17590 -440
rect 6610 -690 17590 -515
rect -800 -815 5785 -770
rect 5820 -710 6580 -700
rect 5820 -770 5830 -710
rect 5980 -770 6420 -710
rect 6570 -770 6580 -710
rect 5820 -780 6580 -770
rect 6610 -770 7220 -690
rect 7580 -770 17590 -690
rect -800 -2375 -780 -815
rect -420 -2375 -380 -815
rect -20 -2375 1220 -815
rect 1580 -2375 5220 -815
rect 5580 -2375 5785 -815
rect -800 -2385 5785 -2375
rect 2005 -2440 2395 -2385
rect 2005 -2515 2025 -2440
rect 2375 -2515 2395 -2440
rect 2005 -2535 2395 -2515
rect 5205 -2440 5595 -2385
rect 5205 -2515 5225 -2440
rect 5575 -2515 5595 -2440
rect 5205 -2535 5595 -2515
rect 2010 -3195 2390 -3180
rect 2010 -3270 2025 -3195
rect 2375 -3270 2390 -3195
rect -800 -3325 830 -3320
rect 2010 -3325 2390 -3270
rect 4410 -3325 4790 -3180
rect 5210 -3195 5590 -3180
rect 5210 -3270 5225 -3195
rect 5575 -3270 5590 -3195
rect 5210 -3325 5590 -3270
rect 6010 -3185 6390 -780
rect 6610 -815 17590 -770
rect 6610 -2375 9220 -815
rect 9580 -2375 10020 -815
rect 10380 -2375 10820 -815
rect 11180 -2375 11220 -815
rect 11580 -2375 11620 -815
rect 11980 -2375 14020 -815
rect 14380 -2375 16420 -815
rect 16780 -2375 16820 -815
rect 17180 -2375 17590 -815
rect 18010 1585 18800 1595
rect 18010 25 18020 1585
rect 18380 25 18420 1585
rect 18780 25 18800 1585
rect 18010 -815 18800 25
rect 18010 -2305 18020 -815
rect 6610 -2385 17590 -2375
rect 18005 -2375 18020 -2305
rect 18380 -2375 18420 -815
rect 18780 -2375 18800 -815
rect 18005 -2385 18800 -2375
rect 19200 1585 19600 1635
rect 19200 25 19220 1585
rect 19580 25 19600 1585
rect 19200 -815 19600 25
rect 19200 -2375 19220 -815
rect 19580 -2375 19600 -815
rect 19200 -2385 19600 -2375
rect 8405 -2440 8795 -2385
rect 8405 -2515 8425 -2440
rect 8775 -2515 8795 -2440
rect 12410 -2515 12790 -2385
rect 14005 -2440 14395 -2385
rect 14005 -2515 14025 -2440
rect 14375 -2515 14395 -2440
rect 15610 -2515 15990 -2385
rect 8405 -2540 8795 -2515
rect 14005 -2540 14395 -2515
rect 6010 -3265 6020 -3185
rect 6380 -3265 6390 -3185
rect 6010 -3275 6390 -3265
rect 6420 -3325 6780 -2740
rect 8410 -3195 8790 -3180
rect 8410 -3270 8425 -3195
rect 8775 -3270 8790 -3195
rect 8410 -3325 8790 -3270
rect 14010 -3190 14390 -3175
rect 14010 -3265 14025 -3190
rect 14375 -3265 14390 -3190
rect 12410 -3325 12790 -3295
rect 14010 -3325 14390 -3265
rect 15610 -3325 15990 -3295
rect 18005 -3325 18790 -2385
rect -800 -3335 18800 -3325
rect -800 -4895 -780 -3335
rect -420 -4895 -380 -3335
rect -20 -4895 4420 -3335
rect 4780 -4895 8420 -3335
rect 8780 -4895 10820 -3335
rect 11180 -4895 11220 -3335
rect 11580 -4895 11620 -3335
rect 11980 -4895 14020 -3335
rect 14380 -4895 16420 -3335
rect 16780 -4895 16820 -3335
rect 17180 -4895 18020 -3335
rect 18380 -4895 18420 -3335
rect 18780 -4895 18800 -3335
rect -800 -4940 18800 -4895
rect 19210 -3335 19600 -2385
rect 19210 -4895 19220 -3335
rect 19580 -4895 19600 -3335
rect 19210 -4905 19600 -4895
rect 20000 1725 20390 1740
rect 20000 1650 20025 1725
rect 20375 1650 20390 1725
rect 20000 5 20390 1650
rect 21600 1725 22000 1740
rect 21600 1650 21625 1725
rect 21975 1650 22000 1725
rect 20800 1585 21195 1605
rect 20800 25 20820 1585
rect 21180 25 21195 1585
rect 20000 -400 20400 5
rect 20000 -475 20025 -400
rect 20375 -475 20400 -400
rect 20000 -2780 20400 -475
rect 20000 -2855 20025 -2780
rect 20375 -2855 20400 -2780
rect -800 -5025 6420 -4940
rect 6780 -5025 18800 -4940
rect -800 -5030 18800 -5025
rect 20000 -5030 20400 -2855
rect -800 -5095 20400 -5030
rect -800 -5140 19280 -5095
rect -800 -5145 4425 -5140
rect -800 -5220 1225 -5145
rect 1575 -5220 4425 -5145
rect -800 -5490 4425 -5220
rect 4775 -5490 6425 -5140
rect 6775 -5490 8425 -5140
rect 8775 -5180 19280 -5140
rect 8775 -5490 14025 -5180
rect -800 -5530 14025 -5490
rect 14375 -5445 19280 -5180
rect 19630 -5165 20400 -5095
rect 20800 -815 21195 25
rect 20800 -2375 20820 -815
rect 21180 -2375 21195 -815
rect 20800 -3335 21195 -2375
rect 20800 -4895 20820 -3335
rect 21180 -4895 21195 -3335
rect 19630 -5445 20405 -5165
rect 14375 -5530 20405 -5445
rect -800 -5605 20405 -5530
rect -800 -5690 6420 -5605
rect 6780 -5690 20405 -5605
rect -800 -5735 20405 -5690
rect -800 -6820 -780 -5735
rect -805 -7295 -780 -6820
rect -420 -7295 -380 -5735
rect -20 -7295 4420 -5735
rect 4780 -7295 8420 -5735
rect 8780 -7295 10820 -5735
rect 11180 -7295 11220 -5735
rect 11580 -7295 11620 -5735
rect 11980 -7295 14015 -5735
rect 14380 -7295 16420 -5735
rect 16780 -7295 16820 -5735
rect 17180 -7295 18020 -5735
rect 18380 -5740 19220 -5735
rect 18380 -7295 18420 -5740
rect -805 -7300 18420 -7295
rect 18780 -7295 19220 -5740
rect 19580 -7295 20405 -5735
rect 18780 -7300 20405 -7295
rect -805 -7360 20405 -7300
rect 20800 -5545 21195 -4895
rect 21600 -385 22000 1650
rect 21600 -460 21635 -385
rect 21985 -460 22000 -385
rect 21600 -2765 22000 -460
rect 22400 1640 24000 1900
rect 22400 1585 22795 1640
rect 22400 25 22420 1585
rect 22780 25 22795 1585
rect 22400 -815 22795 25
rect 22400 -2375 22420 -815
rect 22780 -2375 22795 -815
rect 22400 -2385 22795 -2375
rect 23200 1585 24000 1605
rect 23200 25 23220 1585
rect 23580 25 23620 1585
rect 23980 25 24000 1585
rect 23200 -470 24000 25
rect 23200 -815 24005 -470
rect 23200 -2375 23220 -815
rect 23580 -2375 23620 -815
rect 23980 -2375 24005 -815
rect 23200 -2385 24005 -2375
rect 21600 -2840 21625 -2765
rect 21975 -2840 22000 -2765
rect 21600 -5030 22000 -2840
rect 22410 -3335 22790 -2385
rect 22410 -4895 22420 -3335
rect 22780 -4895 22790 -3335
rect 22410 -4905 22790 -4895
rect 23205 -3335 24005 -2385
rect 23205 -4895 23220 -3335
rect 23580 -4895 23620 -3335
rect 23980 -4895 24005 -3335
rect 23205 -5030 24005 -4895
rect 21600 -5110 24000 -5030
rect 21600 -5460 22340 -5110
rect 22690 -5460 24000 -5110
rect 20800 -5645 21200 -5545
rect 20800 -5735 21195 -5645
rect 20800 -7295 20820 -5735
rect 21180 -7295 21195 -5735
rect 20800 -7315 21195 -7295
rect 21600 -5735 24000 -5460
rect 21600 -7295 22420 -5735
rect 22780 -7295 23220 -5735
rect 23580 -7295 23620 -5735
rect 23980 -7295 24000 -5735
rect 21600 -7305 24000 -7295
rect -805 -7435 2025 -7360
rect 2375 -7435 3625 -7360
rect 3975 -7435 6025 -7360
rect 6375 -7425 8430 -7360
rect 8770 -7425 20405 -7360
rect 6375 -7435 20405 -7425
rect -805 -7455 20405 -7435
rect 20820 -7360 21180 -7350
rect 20820 -7425 20830 -7360
rect 21170 -7425 21180 -7360
rect 20820 -7455 21180 -7425
rect 21610 -7455 24000 -7305
rect -805 -8300 24000 -7455
<< labels >>
rlabel metal1 -805 -7930 -805 -7930 7 GND
rlabel locali -795 -5325 -795 -5325 7 Vr
rlabel metal1 -800 -475 -800 -475 7 VDD
rlabel locali 24000 -7505 24000 -7505 3 Vbn
rlabel locali 23950 -3010 23950 -3010 3 Vg
rlabel metal1 6010 -3010 6010 -3010 7 Vdp
rlabel metal1 21195 -5305 21195 -5305 3 net9
rlabel locali 20995 -655 20995 -655 1 net10
rlabel locali 20990 -3175 20990 -3175 1 net13
rlabel locali 20995 -135 20995 -135 5 net11
rlabel poly 9200 -170 9200 -170 3 Vbp
<< end >>
