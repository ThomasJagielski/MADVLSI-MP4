magic
tech sky130A
magscale 1 2
timestamp 1617054279
<< error_p >>
rect 2353 0 2400 3200
rect 3000 0 3600 3200
rect 4200 0 4800 3200
rect 5400 0 6000 3200
rect 6600 0 7200 3200
rect 7800 0 8400 3200
rect 9000 0 9600 3200
rect 10200 0 10800 3200
rect 11400 0 12000 3200
rect 12600 0 13200 3200
rect 13800 0 14400 3200
rect 15000 0 15600 3200
rect 16200 0 16800 3200
rect 17400 0 18000 3200
rect 18600 0 19200 3200
rect 19800 0 19847 3200
rect 2353 -4000 2400 -800
rect 3000 -4000 3600 -800
rect 4200 -4000 4800 -800
rect 5400 -4000 6000 -800
rect 6600 -4000 7200 -800
rect 7800 -4000 8400 -800
rect 9000 -4000 9600 -800
rect 10200 -4000 10800 -800
rect 11400 -4000 12000 -800
rect 12600 -4000 13200 -800
rect 13800 -4000 14400 -800
rect 15000 -4000 15600 -800
rect 16200 -4000 16800 -800
rect 17400 -4000 18000 -800
rect 18600 -4000 19200 -800
rect 19800 -4000 19847 -800
rect 7800 -8000 8400 -4800
rect 9000 -8000 9600 -4800
rect 10200 -8000 10800 -4800
rect 11400 -8000 12000 -4800
rect 12600 -8000 13200 -4800
rect 13800 -8000 14400 -4800
rect 15000 -8000 15600 -4800
rect 16200 -8000 16800 -4800
rect 17400 -8000 18000 -4800
rect 18600 -8000 19200 -4800
rect 19800 -8000 19847 -4800
<< nmos >>
rect 0 0 600 3200
rect 1200 0 1800 3200
rect 2400 0 3000 3200
rect 3600 0 4200 3200
rect 4800 0 5400 3200
rect 6000 0 6600 3200
rect 7200 0 7800 3200
rect 8400 0 9000 3200
rect 9600 0 10200 3200
rect 10800 0 11400 3200
rect 12000 0 12600 3200
rect 13200 0 13800 3200
rect 14400 0 15000 3200
rect 15600 0 16200 3200
rect 16800 0 17400 3200
rect 18000 0 18600 3200
rect 19200 0 19800 3200
rect 20400 0 21000 3200
rect 21600 0 22200 3200
rect 0 -4000 600 -800
rect 1200 -4000 1800 -800
rect 2400 -4000 3000 -800
rect 3600 -4000 4200 -800
rect 4800 -4000 5400 -800
rect 6000 -4000 6600 -800
rect 7200 -4000 7800 -800
rect 8400 -4000 9000 -800
rect 9600 -4000 10200 -800
rect 10800 -4000 11400 -800
rect 12000 -4000 12600 -800
rect 13200 -4000 13800 -800
rect 14400 -4000 15000 -800
rect 15600 -4000 16200 -800
rect 16800 -4000 17400 -800
rect 18000 -4000 18600 -800
rect 19200 -4000 19800 -800
rect 20400 -4000 21000 -800
rect 21600 -4000 22200 -800
rect 0 -8000 600 -4800
rect 1200 -8000 1800 -4800
rect 2400 -8000 3000 -4800
rect 3600 -8000 4200 -4800
rect 4800 -8000 5400 -4800
rect 6000 -8000 6600 -4800
rect 7200 -8000 7800 -4800
rect 8400 -8000 9000 -4800
rect 9600 -8000 10200 -4800
rect 10800 -8000 11400 -4800
rect 12000 -8000 12600 -4800
rect 13200 -8000 13800 -4800
rect 14400 -8000 15000 -4800
rect 15600 -8000 16200 -4800
rect 16800 -8000 17400 -4800
rect 18000 -8000 18600 -4800
rect 19200 -8000 19800 -4800
rect 20400 -8000 21000 -4800
rect 21600 -8000 22200 -4800
<< ndiff >>
rect -600 3170 0 3200
rect -600 30 -570 3170
rect -30 30 0 3170
rect -600 0 0 30
rect 600 3170 1200 3200
rect 600 30 630 3170
rect 1170 30 1200 3170
rect 600 0 1200 30
rect 1800 3170 2400 3200
rect 1800 30 1830 3170
rect 2370 30 2400 3170
rect 1800 0 2400 30
rect 3000 3170 3600 3200
rect 3000 30 3030 3170
rect 3570 30 3600 3170
rect 3000 0 3600 30
rect 4200 3170 4800 3200
rect 4200 30 4230 3170
rect 4770 30 4800 3170
rect 4200 0 4800 30
rect 5400 3170 6000 3200
rect 5400 30 5430 3170
rect 5970 30 6000 3170
rect 5400 0 6000 30
rect 6600 3170 7200 3200
rect 6600 30 6630 3170
rect 7170 30 7200 3170
rect 6600 0 7200 30
rect 7800 3170 8400 3200
rect 7800 30 7830 3170
rect 8370 30 8400 3170
rect 7800 0 8400 30
rect 9000 3170 9600 3200
rect 9000 30 9030 3170
rect 9570 30 9600 3170
rect 9000 0 9600 30
rect 10200 3170 10800 3200
rect 10200 30 10230 3170
rect 10770 30 10800 3170
rect 10200 0 10800 30
rect 11400 3170 12000 3200
rect 11400 30 11430 3170
rect 11970 30 12000 3170
rect 11400 0 12000 30
rect 12600 3170 13200 3200
rect 12600 30 12630 3170
rect 13170 30 13200 3170
rect 12600 0 13200 30
rect 13800 3170 14400 3200
rect 13800 30 13830 3170
rect 14370 30 14400 3170
rect 13800 0 14400 30
rect 15000 3170 15600 3200
rect 15000 30 15030 3170
rect 15570 30 15600 3170
rect 15000 0 15600 30
rect 16200 3170 16800 3200
rect 16200 30 16230 3170
rect 16770 30 16800 3170
rect 16200 0 16800 30
rect 17400 3170 18000 3200
rect 17400 30 17430 3170
rect 17970 30 18000 3170
rect 17400 0 18000 30
rect 18600 3170 19200 3200
rect 18600 30 18630 3170
rect 19170 30 19200 3170
rect 18600 0 19200 30
rect 19800 3170 20400 3200
rect 19800 30 19830 3170
rect 20370 30 20400 3170
rect 19800 0 20400 30
rect 21000 3170 21600 3200
rect 21000 30 21030 3170
rect 21570 30 21600 3170
rect 21000 0 21600 30
rect 22200 3170 22800 3200
rect 22200 30 22230 3170
rect 22770 30 22800 3170
rect 22200 0 22800 30
rect -600 -830 0 -800
rect -600 -3970 -570 -830
rect -30 -3970 0 -830
rect -600 -4000 0 -3970
rect 600 -830 1200 -800
rect 600 -3970 630 -830
rect 1170 -3970 1200 -830
rect 600 -4000 1200 -3970
rect 1800 -830 2400 -800
rect 1800 -3970 1830 -830
rect 2370 -3970 2400 -830
rect 1800 -4000 2400 -3970
rect 3000 -830 3600 -800
rect 3000 -3970 3030 -830
rect 3570 -3970 3600 -830
rect 3000 -4000 3600 -3970
rect 4200 -830 4800 -800
rect 4200 -3970 4230 -830
rect 4770 -3970 4800 -830
rect 4200 -4000 4800 -3970
rect 5400 -830 6000 -800
rect 5400 -3970 5430 -830
rect 5970 -3970 6000 -830
rect 5400 -4000 6000 -3970
rect 6600 -830 7200 -800
rect 6600 -3970 6630 -830
rect 7170 -3970 7200 -830
rect 6600 -4000 7200 -3970
rect 7800 -830 8400 -800
rect 7800 -3970 7830 -830
rect 8370 -3970 8400 -830
rect 7800 -4000 8400 -3970
rect 9000 -830 9600 -800
rect 9000 -3970 9030 -830
rect 9570 -3970 9600 -830
rect 9000 -4000 9600 -3970
rect 10200 -830 10800 -800
rect 10200 -3970 10230 -830
rect 10770 -3970 10800 -830
rect 10200 -4000 10800 -3970
rect 11400 -830 12000 -800
rect 11400 -3970 11430 -830
rect 11970 -3970 12000 -830
rect 11400 -4000 12000 -3970
rect 12600 -830 13200 -800
rect 12600 -3970 12630 -830
rect 13170 -3970 13200 -830
rect 12600 -4000 13200 -3970
rect 13800 -830 14400 -800
rect 13800 -3970 13830 -830
rect 14370 -3970 14400 -830
rect 13800 -4000 14400 -3970
rect 15000 -830 15600 -800
rect 15000 -3970 15030 -830
rect 15570 -3970 15600 -830
rect 15000 -4000 15600 -3970
rect 16200 -830 16800 -800
rect 16200 -3970 16230 -830
rect 16770 -3970 16800 -830
rect 16200 -4000 16800 -3970
rect 17400 -830 18000 -800
rect 17400 -3970 17430 -830
rect 17970 -3970 18000 -830
rect 17400 -4000 18000 -3970
rect 18600 -830 19200 -800
rect 18600 -3970 18630 -830
rect 19170 -3970 19200 -830
rect 18600 -4000 19200 -3970
rect 19800 -830 20400 -800
rect 19800 -3970 19830 -830
rect 20370 -3970 20400 -830
rect 19800 -4000 20400 -3970
rect 21000 -830 21600 -800
rect 21000 -3970 21030 -830
rect 21570 -3970 21600 -830
rect 21000 -4000 21600 -3970
rect 22200 -830 22800 -800
rect 22200 -3970 22230 -830
rect 22770 -3970 22800 -830
rect 22200 -4000 22800 -3970
rect -600 -4830 0 -4800
rect -600 -7970 -570 -4830
rect -30 -7970 0 -4830
rect -600 -8000 0 -7970
rect 600 -4830 1200 -4800
rect 600 -7970 630 -4830
rect 1170 -7970 1200 -4830
rect 600 -8000 1200 -7970
rect 1800 -4830 2400 -4800
rect 1800 -7970 1830 -4830
rect 2370 -7970 2400 -4830
rect 1800 -8000 2400 -7970
rect 3000 -4830 3600 -4800
rect 3000 -7970 3030 -4830
rect 3570 -7970 3600 -4830
rect 3000 -8000 3600 -7970
rect 4200 -4830 4800 -4800
rect 4200 -7970 4230 -4830
rect 4770 -7970 4800 -4830
rect 4200 -8000 4800 -7970
rect 5400 -4830 6000 -4800
rect 5400 -7970 5430 -4830
rect 5970 -7970 6000 -4830
rect 5400 -8000 6000 -7970
rect 6600 -4830 7200 -4800
rect 6600 -7970 6630 -4830
rect 7170 -7970 7200 -4830
rect 6600 -8000 7200 -7970
rect 7800 -4830 8400 -4800
rect 7800 -7970 7830 -4830
rect 8370 -7970 8400 -4830
rect 7800 -8000 8400 -7970
rect 9000 -4830 9600 -4800
rect 9000 -7970 9030 -4830
rect 9570 -7970 9600 -4830
rect 9000 -8000 9600 -7970
rect 10200 -4830 10800 -4800
rect 10200 -7970 10230 -4830
rect 10770 -7970 10800 -4830
rect 10200 -8000 10800 -7970
rect 11400 -4830 12000 -4800
rect 11400 -7970 11430 -4830
rect 11970 -7970 12000 -4830
rect 11400 -8000 12000 -7970
rect 12600 -4830 13200 -4800
rect 12600 -7970 12630 -4830
rect 13170 -7970 13200 -4830
rect 12600 -8000 13200 -7970
rect 13800 -4830 14400 -4800
rect 13800 -7970 13830 -4830
rect 14370 -7970 14400 -4830
rect 13800 -8000 14400 -7970
rect 15000 -4830 15600 -4800
rect 15000 -7970 15030 -4830
rect 15570 -7970 15600 -4830
rect 15000 -8000 15600 -7970
rect 16200 -4830 16800 -4800
rect 16200 -7970 16230 -4830
rect 16770 -7970 16800 -4830
rect 16200 -8000 16800 -7970
rect 17400 -4830 18000 -4800
rect 17400 -7970 17430 -4830
rect 17970 -7970 18000 -4830
rect 17400 -8000 18000 -7970
rect 18600 -4830 19200 -4800
rect 18600 -7970 18630 -4830
rect 19170 -7970 19200 -4830
rect 18600 -8000 19200 -7970
rect 19800 -4830 20400 -4800
rect 19800 -7970 19830 -4830
rect 20370 -7970 20400 -4830
rect 19800 -8000 20400 -7970
rect 21000 -4830 21600 -4800
rect 21000 -7970 21030 -4830
rect 21570 -7970 21600 -4830
rect 21000 -8000 21600 -7970
rect 22200 -4830 22800 -4800
rect 22200 -7970 22230 -4830
rect 22770 -7970 22800 -4830
rect 22200 -8000 22800 -7970
<< ndiffc >>
rect -570 30 -30 3170
rect 630 30 1170 3170
rect 1830 30 2370 3170
rect 3030 30 3570 3170
rect 4230 30 4770 3170
rect 5430 30 5970 3170
rect 6630 30 7170 3170
rect 7830 30 8370 3170
rect 9030 30 9570 3170
rect 10230 30 10770 3170
rect 11430 30 11970 3170
rect 12630 30 13170 3170
rect 13830 30 14370 3170
rect 15030 30 15570 3170
rect 16230 30 16770 3170
rect 17430 30 17970 3170
rect 18630 30 19170 3170
rect 19830 30 20370 3170
rect 21030 30 21570 3170
rect 22230 30 22770 3170
rect -570 -3970 -30 -830
rect 630 -3970 1170 -830
rect 1830 -3970 2370 -830
rect 3030 -3970 3570 -830
rect 4230 -3970 4770 -830
rect 5430 -3970 5970 -830
rect 6630 -3970 7170 -830
rect 7830 -3970 8370 -830
rect 9030 -3970 9570 -830
rect 10230 -3970 10770 -830
rect 11430 -3970 11970 -830
rect 12630 -3970 13170 -830
rect 13830 -3970 14370 -830
rect 15030 -3970 15570 -830
rect 16230 -3970 16770 -830
rect 17430 -3970 17970 -830
rect 18630 -3970 19170 -830
rect 19830 -3970 20370 -830
rect 21030 -3970 21570 -830
rect 22230 -3970 22770 -830
rect -570 -7970 -30 -4830
rect 630 -7970 1170 -4830
rect 1830 -7970 2370 -4830
rect 3030 -7970 3570 -4830
rect 4230 -7970 4770 -4830
rect 5430 -7970 5970 -4830
rect 6630 -7970 7170 -4830
rect 7830 -7970 8370 -4830
rect 9030 -7970 9570 -4830
rect 10230 -7970 10770 -4830
rect 11430 -7970 11970 -4830
rect 12630 -7970 13170 -4830
rect 13830 -7970 14370 -4830
rect 15030 -7970 15570 -4830
rect 16230 -7970 16770 -4830
rect 17430 -7970 17970 -4830
rect 18630 -7970 19170 -4830
rect 19830 -7970 20370 -4830
rect 21030 -7970 21570 -4830
rect 22230 -7970 22770 -4830
<< psubdiff >>
rect -1200 3170 -600 3200
rect -1200 30 -1170 3170
rect -630 30 -600 3170
rect -1200 0 -600 30
rect 22800 3170 23400 3200
rect 22800 30 22830 3170
rect 23370 30 23400 3170
rect 22800 0 23400 30
rect -1200 -830 -600 -800
rect -1200 -3970 -1170 -830
rect -630 -3970 -600 -830
rect -1200 -4000 -600 -3970
rect 22800 -830 23400 -800
rect 22800 -3970 22830 -830
rect 23370 -3970 23400 -830
rect 22800 -4000 23400 -3970
rect -1200 -4830 -600 -4800
rect -1200 -7970 -1170 -4830
rect -630 -7970 -600 -4830
rect -1200 -8000 -600 -7970
rect 22800 -4830 23400 -4800
rect 22800 -7970 22830 -4830
rect 23370 -7970 23400 -4830
rect 22800 -8000 23400 -7970
<< psubdiffcont >>
rect -1170 30 -630 3170
rect 22830 30 23370 3170
rect -1170 -3970 -630 -830
rect 22830 -3970 23370 -830
rect -1170 -7970 -630 -4830
rect 22830 -7970 23370 -4830
<< poly >>
rect 860 3290 940 3310
rect 860 3260 880 3290
rect 0 3250 880 3260
rect 920 3260 940 3290
rect 2400 3280 19800 3310
rect 920 3250 1800 3260
rect 0 3230 1800 3250
rect 0 3200 600 3230
rect 1200 3200 1800 3230
rect 2400 3200 3000 3280
rect 3600 3200 4200 3280
rect 4800 3200 5400 3230
rect 6000 3200 6600 3280
rect 7200 3200 7800 3230
rect 8400 3200 9000 3280
rect 9600 3200 10200 3230
rect 10800 3200 11400 3280
rect 12000 3200 12600 3230
rect 13200 3200 13800 3280
rect 14400 3200 15000 3230
rect 15600 3200 16200 3280
rect 16800 3200 17400 3230
rect 18000 3200 18600 3280
rect 19200 3200 19800 3280
rect 21240 3290 21320 3310
rect 21240 3260 21260 3290
rect 20400 3250 21260 3260
rect 21300 3260 21320 3290
rect 21300 3250 22200 3260
rect 20400 3230 22200 3250
rect 20400 3200 21000 3230
rect 21600 3200 22200 3230
rect 0 -30 600 0
rect 1200 -30 1800 0
rect 2400 -30 3000 0
rect 3600 -30 4200 0
rect 4800 -30 5400 0
rect 6000 -30 6600 0
rect 7200 -30 7800 0
rect 8400 -30 9000 0
rect 9600 -30 10200 0
rect 10800 -30 11400 0
rect 12000 -30 12600 0
rect 13200 -30 13800 0
rect 14400 -30 15000 0
rect 15600 -30 16200 0
rect 16800 -30 17400 0
rect 18000 -30 18600 0
rect 19200 -30 19800 0
rect 20400 -30 21000 0
rect 21600 -30 22200 0
rect 0 -800 600 -770
rect 1200 -800 1800 -770
rect 2400 -800 3000 -770
rect 3600 -800 4200 -770
rect 4800 -800 5400 -770
rect 6000 -800 6600 -770
rect 7200 -800 7800 -770
rect 8400 -800 9000 -770
rect 9600 -800 10200 -770
rect 10800 -800 11400 -770
rect 12000 -800 12600 -770
rect 13200 -800 13800 -770
rect 14400 -800 15000 -770
rect 15600 -800 16200 -770
rect 16800 -800 17400 -770
rect 18000 -800 18600 -770
rect 19200 -800 19800 -770
rect 20400 -800 21000 -770
rect 21600 -800 22200 -770
rect 0 -4030 600 -4000
rect 1200 -4030 1800 -4000
rect 2400 -4030 3000 -4000
rect 3600 -4030 4200 -4000
rect 4800 -4030 5400 -4000
rect 6000 -4030 6600 -4000
rect 7200 -4030 7800 -4000
rect 8400 -4030 9000 -4000
rect 9600 -4030 10200 -4000
rect 10800 -4030 11400 -4000
rect 12000 -4030 12600 -4000
rect 13200 -4030 13800 -4000
rect 14400 -4030 15000 -4000
rect 15600 -4030 16200 -4000
rect 16800 -4030 17400 -4000
rect 18000 -4030 18600 -4000
rect 19200 -4030 19800 -4000
rect 20400 -4030 21000 -4000
rect 21600 -4030 22200 -4000
rect 0 -4800 600 -4770
rect 1200 -4800 1800 -4770
rect 2400 -4800 3000 -4770
rect 3600 -4800 4200 -4770
rect 4800 -4800 5400 -4770
rect 6000 -4800 6600 -4770
rect 7200 -4800 7800 -4770
rect 8400 -4800 9000 -4770
rect 9600 -4800 10200 -4770
rect 10800 -4800 11400 -4770
rect 12000 -4800 12600 -4770
rect 13200 -4800 13800 -4770
rect 14400 -4800 15000 -4770
rect 15600 -4800 16200 -4770
rect 16800 -4800 17400 -4770
rect 18000 -4800 18600 -4770
rect 19200 -4800 19800 -4770
rect 20400 -4800 21000 -4770
rect 21600 -4800 22200 -4770
rect 0 -8030 600 -8000
rect 1200 -8030 1800 -8000
rect 2400 -8030 3000 -8000
rect 3600 -8030 4200 -8000
rect 4800 -8030 5400 -8000
rect 6000 -8030 6600 -8000
rect 7200 -8030 7800 -8000
rect 8400 -8030 9000 -8000
rect 9600 -8030 10200 -8000
rect 10800 -8030 11400 -8000
rect 12000 -8030 12600 -8000
rect 13200 -8030 13800 -8000
rect 14400 -8030 15000 -8000
rect 15600 -8030 16200 -8000
rect 16800 -8030 17400 -8000
rect 18000 -8030 18600 -8000
rect 19200 -8030 19800 -8000
rect 20400 -8030 21000 -8000
rect 21600 -8030 22200 -8000
<< polycont >>
rect 880 3250 920 3290
rect 21260 3250 21300 3290
<< locali >>
rect 18610 3360 23400 3400
rect 860 3290 940 3310
rect 860 3250 880 3290
rect 920 3250 940 3290
rect 860 3230 940 3250
rect -1190 3170 -10 3190
rect -1190 30 -1170 3170
rect -630 30 -570 3170
rect -30 30 -10 3170
rect -1190 10 -10 30
rect 610 3170 1190 3230
rect 610 30 630 3170
rect 1170 30 1190 3170
rect 610 10 1190 30
rect 1810 3170 2390 3190
rect 1810 30 1830 3170
rect 2370 30 2390 3170
rect 1810 -40 2390 30
rect 3010 3170 3590 3190
rect 3010 30 3030 3170
rect 3570 30 3590 3170
rect 3010 10 3590 30
rect 4210 3170 4790 3190
rect 4210 30 4230 3170
rect 4770 30 4790 3170
rect 4210 -40 4790 30
rect 1810 -80 4790 -40
rect 5410 3170 5990 3190
rect 5410 30 5430 3170
rect 5970 30 5990 3170
rect 5410 -80 5990 30
rect 6610 3170 7190 3190
rect 6610 30 6630 3170
rect 7170 30 7190 3170
rect 6610 10 7190 30
rect 7810 3170 8390 3190
rect 7810 30 7830 3170
rect 8370 30 8390 3170
rect 7810 10 8390 30
rect 9010 3170 9590 3190
rect 9010 30 9030 3170
rect 9570 30 9590 3170
rect 9010 -80 9590 30
rect 10210 3170 10790 3190
rect 10210 30 10230 3170
rect 10770 30 10790 3170
rect 10210 -70 10790 30
rect 11410 3170 11990 3190
rect 11410 30 11430 3170
rect 11970 30 11990 3170
rect 11410 10 11990 30
rect 12610 3170 13190 3190
rect 12610 30 12630 3170
rect 13170 30 13190 3170
rect 12610 -70 13190 30
rect 13810 3170 14390 3190
rect 13810 30 13830 3170
rect 14370 30 14390 3170
rect 13810 10 14390 30
rect 15010 3170 15590 3190
rect 15010 30 15030 3170
rect 15570 30 15590 3170
rect 15010 -70 15590 30
rect 16210 3170 16790 3190
rect 16210 30 16230 3170
rect 16770 30 16790 3170
rect 16210 10 16790 30
rect 17410 3170 17990 3190
rect 17410 30 17430 3170
rect 17970 30 17990 3170
rect 17410 -40 17990 30
rect 18610 3170 19190 3360
rect 21240 3290 21320 3310
rect 21240 3250 21260 3290
rect 21300 3250 21320 3290
rect 21240 3230 21320 3250
rect 18610 30 18630 3170
rect 19170 30 19190 3170
rect 18610 10 19190 30
rect 19810 3170 20390 3190
rect 19810 30 19830 3170
rect 20370 30 20390 3170
rect 19810 -40 20390 30
rect 21010 3170 21590 3230
rect 21010 30 21030 3170
rect 21570 30 21590 3170
rect 21010 10 21590 30
rect 22210 3170 23390 3190
rect 22210 30 22230 3170
rect 22770 30 22830 3170
rect 23370 30 23390 3170
rect 22210 10 23390 30
rect 3300 -270 3340 -80
rect 5680 -210 5720 -80
rect 9280 -250 9320 -80
rect 10480 -250 10520 -70
rect 12880 -250 12920 -70
rect 15280 -250 15320 -70
rect 17410 -80 20390 -40
rect 18890 -310 18930 -80
rect -1190 -830 -10 -810
rect -1190 -3970 -1170 -830
rect -630 -3970 -570 -830
rect -30 -3970 -10 -830
rect -1190 -3990 -10 -3970
rect 610 -830 1190 -810
rect 610 -3970 630 -830
rect 1170 -3970 1190 -830
rect 610 -3990 1190 -3970
rect 1810 -830 2390 -810
rect 1810 -3970 1830 -830
rect 2370 -3970 2390 -830
rect 1810 -3990 2390 -3970
rect 3010 -830 3590 -810
rect 3010 -3970 3030 -830
rect 3570 -3970 3590 -830
rect 3010 -3990 3590 -3970
rect 4210 -830 4790 -810
rect 4210 -3970 4230 -830
rect 4770 -3970 4790 -830
rect 4210 -3990 4790 -3970
rect 5410 -830 5990 -810
rect 5410 -3970 5430 -830
rect 5970 -3970 5990 -830
rect 5410 -3990 5990 -3970
rect 6610 -830 7190 -810
rect 6610 -3970 6630 -830
rect 7170 -3970 7190 -830
rect 6610 -3990 7190 -3970
rect 7810 -830 8390 -810
rect 7810 -3970 7830 -830
rect 8370 -3970 8390 -830
rect 7810 -3990 8390 -3970
rect 9010 -830 9590 -810
rect 9010 -3970 9030 -830
rect 9570 -3970 9590 -830
rect 9010 -3990 9590 -3970
rect 10210 -830 10790 -810
rect 10210 -3970 10230 -830
rect 10770 -3970 10790 -830
rect 10210 -3990 10790 -3970
rect 11410 -830 11990 -810
rect 11410 -3970 11430 -830
rect 11970 -3970 11990 -830
rect 11410 -3990 11990 -3970
rect 12610 -830 13190 -810
rect 12610 -3970 12630 -830
rect 13170 -3970 13190 -830
rect 12610 -3990 13190 -3970
rect 13810 -830 14390 -810
rect 13810 -3970 13830 -830
rect 14370 -3970 14390 -830
rect 13810 -3990 14390 -3970
rect 15010 -830 15590 -810
rect 15010 -3970 15030 -830
rect 15570 -3970 15590 -830
rect 15010 -3990 15590 -3970
rect 16210 -830 16790 -810
rect 16210 -3970 16230 -830
rect 16770 -3970 16790 -830
rect 16210 -3990 16790 -3970
rect 17410 -830 17990 -810
rect 17410 -3970 17430 -830
rect 17970 -3970 17990 -830
rect 17410 -3990 17990 -3970
rect 18610 -830 19190 -810
rect 18610 -3970 18630 -830
rect 19170 -3970 19190 -830
rect 18610 -3990 19190 -3970
rect 19810 -830 20390 -810
rect 19810 -3970 19830 -830
rect 20370 -3970 20390 -830
rect 19810 -3990 20390 -3970
rect 21010 -830 21590 -810
rect 21010 -3970 21030 -830
rect 21570 -3970 21590 -830
rect 21010 -3990 21590 -3970
rect 22210 -830 23390 -810
rect 22210 -3970 22230 -830
rect 22770 -3970 22830 -830
rect 23370 -3970 23390 -830
rect 22210 -3990 23390 -3970
rect -1190 -4830 -10 -4810
rect -1190 -7970 -1170 -4830
rect -630 -7970 -570 -4830
rect -30 -7970 -10 -4830
rect -1190 -7990 -10 -7970
rect 610 -4830 1190 -4810
rect 610 -7970 630 -4830
rect 1170 -7970 1190 -4830
rect 610 -7990 1190 -7970
rect 1810 -4830 2390 -4810
rect 1810 -7970 1830 -4830
rect 2370 -7970 2390 -4830
rect 1810 -7990 2390 -7970
rect 3010 -4830 3590 -4810
rect 3010 -7970 3030 -4830
rect 3570 -7970 3590 -4830
rect 3010 -7990 3590 -7970
rect 4210 -4830 4790 -4810
rect 4210 -7970 4230 -4830
rect 4770 -7970 4790 -4830
rect 4210 -7990 4790 -7970
rect 5410 -4830 5990 -4810
rect 5410 -7970 5430 -4830
rect 5970 -7970 5990 -4830
rect 5410 -7990 5990 -7970
rect 6610 -4830 7190 -4810
rect 6610 -7970 6630 -4830
rect 7170 -7970 7190 -4830
rect 6610 -7990 7190 -7970
rect 7810 -4830 8390 -4810
rect 7810 -7970 7830 -4830
rect 8370 -7970 8390 -4830
rect 7810 -7990 8390 -7970
rect 9010 -4830 9590 -4810
rect 9010 -7970 9030 -4830
rect 9570 -7970 9590 -4830
rect 9010 -7990 9590 -7970
rect 10210 -4830 10790 -4810
rect 10210 -7970 10230 -4830
rect 10770 -7970 10790 -4830
rect 10210 -7990 10790 -7970
rect 11410 -4830 11990 -4810
rect 11410 -7970 11430 -4830
rect 11970 -7970 11990 -4830
rect 11410 -7990 11990 -7970
rect 12610 -4830 13190 -4810
rect 12610 -7970 12630 -4830
rect 13170 -7970 13190 -4830
rect 12610 -7990 13190 -7970
rect 13810 -4830 14390 -4810
rect 13810 -7970 13830 -4830
rect 14370 -7970 14390 -4830
rect 13810 -7990 14390 -7970
rect 15010 -4830 15590 -4810
rect 15010 -7970 15030 -4830
rect 15570 -7970 15590 -4830
rect 15010 -7990 15590 -7970
rect 16210 -4830 16790 -4810
rect 16210 -7970 16230 -4830
rect 16770 -7970 16790 -4830
rect 16210 -7990 16790 -7970
rect 17410 -4830 17990 -4810
rect 17410 -7970 17430 -4830
rect 17970 -7970 17990 -4830
rect 17410 -7990 17990 -7970
rect 18610 -4830 19190 -4810
rect 18610 -7970 18630 -4830
rect 19170 -7970 19190 -4830
rect 18610 -7990 19190 -7970
rect 19810 -4830 20390 -4810
rect 19810 -7970 19830 -4830
rect 20370 -7970 20390 -4830
rect 19810 -7990 20390 -7970
rect 21010 -4830 21590 -4810
rect 21010 -7970 21030 -4830
rect 21570 -7970 21590 -4830
rect 21010 -7990 21590 -7970
rect 22210 -4830 23390 -4810
rect 22210 -7970 22230 -4830
rect 22770 -7970 22830 -4830
rect 23370 -7970 23390 -4830
rect 22210 -7990 23390 -7970
<< end >>
