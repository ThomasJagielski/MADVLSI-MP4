magic
tech sky130A
magscale 1 2
timestamp 1617104566
<< error_p >>
rect 2353 0 2400 3200
rect 3000 0 3600 3200
rect 4200 0 4800 3200
rect 5400 0 6000 3200
rect 6600 0 7200 3200
rect 7800 0 8400 3200
rect 9000 0 9600 3200
rect 10200 0 10800 3200
rect 11400 0 12000 3200
rect 12600 0 13200 3200
rect 13800 0 14400 3200
rect 15000 0 15600 3200
rect 16200 0 16800 3200
rect 17400 0 18000 3200
rect 18600 0 19200 3200
rect 19800 0 19847 3200
<< nwell >>
rect -1240 -50 23440 3240
<< pmos >>
rect 0 0 600 3200
rect 1200 0 1800 3200
rect 2400 0 3000 3200
rect 3600 0 4200 3200
rect 4800 0 5400 3200
rect 6000 0 6600 3200
rect 7200 0 7800 3200
rect 8400 0 9000 3200
rect 9600 0 10200 3200
rect 10800 0 11400 3200
rect 12000 0 12600 3200
rect 13200 0 13800 3200
rect 14400 0 15000 3200
rect 15600 0 16200 3200
rect 16800 0 17400 3200
rect 18000 0 18600 3200
rect 19200 0 19800 3200
rect 20400 0 21000 3200
rect 21600 0 22200 3200
<< pdiff >>
rect -600 3170 0 3200
rect -600 30 -570 3170
rect -30 30 0 3170
rect -600 0 0 30
rect 600 3170 1200 3200
rect 600 30 630 3170
rect 1170 30 1200 3170
rect 600 0 1200 30
rect 1800 3170 2400 3200
rect 1800 30 1830 3170
rect 2370 30 2400 3170
rect 1800 0 2400 30
rect 3000 3170 3600 3200
rect 3000 30 3030 3170
rect 3570 30 3600 3170
rect 3000 0 3600 30
rect 4200 3170 4800 3200
rect 4200 30 4230 3170
rect 4770 30 4800 3170
rect 4200 0 4800 30
rect 5400 3170 6000 3200
rect 5400 30 5430 3170
rect 5970 30 6000 3170
rect 5400 0 6000 30
rect 6600 3170 7200 3200
rect 6600 30 6630 3170
rect 7170 30 7200 3170
rect 6600 0 7200 30
rect 7800 3170 8400 3200
rect 7800 30 7830 3170
rect 8370 30 8400 3170
rect 7800 0 8400 30
rect 9000 3170 9600 3200
rect 9000 30 9030 3170
rect 9570 30 9600 3170
rect 9000 0 9600 30
rect 10200 3170 10800 3200
rect 10200 30 10230 3170
rect 10770 30 10800 3170
rect 10200 0 10800 30
rect 11400 3170 12000 3200
rect 11400 30 11430 3170
rect 11970 30 12000 3170
rect 11400 0 12000 30
rect 12600 3170 13200 3200
rect 12600 30 12630 3170
rect 13170 30 13200 3170
rect 12600 0 13200 30
rect 13800 3170 14400 3200
rect 13800 30 13830 3170
rect 14370 30 14400 3170
rect 13800 0 14400 30
rect 15000 3170 15600 3200
rect 15000 30 15030 3170
rect 15570 30 15600 3170
rect 15000 0 15600 30
rect 16200 3170 16800 3200
rect 16200 30 16230 3170
rect 16770 30 16800 3170
rect 16200 0 16800 30
rect 17400 3170 18000 3200
rect 17400 30 17430 3170
rect 17970 30 18000 3170
rect 17400 0 18000 30
rect 18600 3170 19200 3200
rect 18600 30 18630 3170
rect 19170 30 19200 3170
rect 18600 0 19200 30
rect 19800 3170 20400 3200
rect 19800 30 19830 3170
rect 20370 30 20400 3170
rect 19800 0 20400 30
rect 21000 3170 21600 3200
rect 21000 30 21030 3170
rect 21570 30 21600 3170
rect 21000 0 21600 30
rect 22200 3170 22800 3200
rect 22200 30 22230 3170
rect 22770 30 22800 3170
rect 22200 0 22800 30
<< pdiffc >>
rect -570 30 -30 3170
rect 630 30 1170 3170
rect 1830 30 2370 3170
rect 3030 30 3570 3170
rect 4230 30 4770 3170
rect 5430 30 5970 3170
rect 6630 30 7170 3170
rect 7830 30 8370 3170
rect 9030 30 9570 3170
rect 10230 30 10770 3170
rect 11430 30 11970 3170
rect 12630 30 13170 3170
rect 13830 30 14370 3170
rect 15030 30 15570 3170
rect 16230 30 16770 3170
rect 17430 30 17970 3170
rect 18630 30 19170 3170
rect 19830 30 20370 3170
rect 21030 30 21570 3170
rect 22230 30 22770 3170
<< nsubdiff >>
rect -1200 3170 -600 3200
rect -1200 30 -1170 3170
rect -630 30 -600 3170
rect -1200 0 -600 30
rect 22800 3170 23400 3200
rect 22800 30 22830 3170
rect 23370 30 23400 3170
rect 22800 0 23400 30
<< nsubdiffcont >>
rect -1170 30 -630 3170
rect 22830 30 23370 3170
<< poly >>
rect -340 3290 -260 3310
rect -340 3260 -320 3290
rect -590 3250 -320 3260
rect -280 3260 -260 3290
rect 860 3290 940 3310
rect 860 3260 880 3290
rect -280 3250 880 3260
rect 920 3260 940 3290
rect 2060 3290 2140 3310
rect 2060 3260 2080 3290
rect 920 3250 2080 3260
rect 2120 3260 2140 3290
rect 3260 3290 3340 3310
rect 3260 3260 3280 3290
rect 2120 3250 3280 3260
rect 3320 3260 3340 3290
rect 20040 3290 20120 3310
rect 20040 3260 20060 3290
rect 3320 3250 4200 3260
rect -590 3230 4200 3250
rect 19200 3250 20060 3260
rect 20100 3260 20120 3290
rect 21240 3290 21320 3310
rect 21240 3260 21260 3290
rect 20100 3250 21260 3260
rect 21300 3260 21320 3290
rect 22460 3290 22540 3310
rect 22460 3260 22480 3290
rect 21300 3250 22480 3260
rect 22520 3260 22540 3290
rect 22520 3250 22790 3260
rect 19200 3230 22790 3250
rect 0 3200 600 3230
rect 1200 3200 1800 3230
rect 2400 3200 3000 3230
rect 3600 3200 4200 3230
rect 4800 3200 5400 3230
rect 6000 3200 6600 3230
rect 7200 3200 7800 3230
rect 8400 3200 9000 3230
rect 9600 3200 10200 3230
rect 10800 3200 11400 3230
rect 12000 3200 12600 3230
rect 13200 3200 13800 3230
rect 14400 3200 15000 3230
rect 15600 3200 16200 3230
rect 16800 3200 17400 3230
rect 18000 3200 18600 3230
rect 19200 3200 19800 3230
rect 20400 3200 21000 3230
rect 21600 3200 22200 3230
rect 0 -30 600 0
rect 1200 -30 1800 0
rect 2400 -30 3000 0
rect 3600 -30 4200 0
rect 4800 -30 5400 0
rect 6000 -30 6600 0
rect 7200 -30 7800 0
rect 8400 -30 9000 0
rect 9600 -30 10200 0
rect 10800 -30 11400 0
rect 12000 -30 12600 0
rect 13200 -30 13800 0
rect 14400 -30 15000 0
rect 15600 -30 16200 0
rect 16800 -30 17400 0
rect 18000 -30 18600 0
rect 19200 -30 19800 0
rect 20400 -30 21000 0
rect 21600 -30 22200 0
<< polycont >>
rect -320 3250 -280 3290
rect 880 3250 920 3290
rect 2080 3250 2120 3290
rect 3280 3250 3320 3290
rect 20060 3250 20100 3290
rect 21260 3250 21300 3290
rect 22480 3250 22520 3290
<< locali >>
rect 4210 3330 19190 3370
rect -340 3290 -260 3310
rect -340 3250 -320 3290
rect -280 3250 -260 3290
rect -340 3230 -260 3250
rect 860 3290 940 3310
rect 860 3250 880 3290
rect 920 3250 940 3290
rect 860 3230 940 3250
rect 2060 3290 2140 3310
rect 2060 3250 2080 3290
rect 2120 3250 2140 3290
rect 2060 3230 2140 3250
rect 3260 3290 3340 3310
rect 3260 3250 3280 3290
rect 3320 3250 3340 3290
rect 3260 3230 3340 3250
rect -590 3190 -10 3230
rect -1190 3170 -10 3190
rect -1190 30 -1170 3170
rect -630 30 -570 3170
rect -30 30 -10 3170
rect -1190 10 -10 30
rect 610 3170 1190 3230
rect 610 30 630 3170
rect 1170 30 1190 3170
rect 610 10 1190 30
rect 1810 3170 2390 3230
rect 1810 30 1830 3170
rect 2370 30 2390 3170
rect 1810 0 2390 30
rect 3010 3170 3590 3230
rect 3010 30 3030 3170
rect 3570 30 3590 3170
rect 3010 10 3590 30
rect 4210 3170 4790 3330
rect 4210 30 4230 3170
rect 4770 30 4790 3170
rect 4210 0 4790 30
rect 5410 3240 17990 3280
rect 5410 3170 5990 3240
rect 5410 30 5430 3170
rect 5970 30 5990 3170
rect 5410 0 5990 30
rect 6610 3170 7190 3190
rect 6610 30 6630 3170
rect 7170 30 7190 3170
rect 6610 10 7190 30
rect 7810 3170 8390 3190
rect 7810 30 7830 3170
rect 8370 30 8390 3170
rect 7810 10 8390 30
rect 9010 3170 9590 3190
rect 9010 30 9030 3170
rect 9570 30 9590 3170
rect 9010 0 9590 30
rect 10210 3170 10790 3240
rect 10210 30 10230 3170
rect 10770 30 10790 3170
rect 10210 0 10790 30
rect 11410 3170 11990 3190
rect 11410 30 11430 3170
rect 11970 30 11990 3170
rect 11410 10 11990 30
rect 12610 3170 13190 3240
rect 12610 30 12630 3170
rect 13170 30 13190 3170
rect 12610 0 13190 30
rect 13810 3170 14390 3190
rect 13810 30 13830 3170
rect 14370 30 14390 3170
rect 13810 10 14390 30
rect 15010 3170 15590 3190
rect 15010 30 15030 3170
rect 15570 30 15590 3170
rect 15010 0 15590 30
rect 16210 3170 16790 3190
rect 16210 30 16230 3170
rect 16770 30 16790 3170
rect 16210 10 16790 30
rect 17410 3170 17990 3240
rect 17410 30 17430 3170
rect 17970 30 17990 3170
rect 17410 0 17990 30
rect 18610 3170 19190 3330
rect 20040 3290 20120 3310
rect 20040 3250 20060 3290
rect 20100 3250 20120 3290
rect 20040 3230 20120 3250
rect 21240 3290 21320 3310
rect 21240 3250 21260 3290
rect 21300 3250 21320 3290
rect 21240 3230 21320 3250
rect 22460 3290 22540 3310
rect 22460 3250 22480 3290
rect 22520 3250 22540 3290
rect 22460 3230 22540 3250
rect 18610 30 18630 3170
rect 19170 30 19190 3170
rect 18610 10 19190 30
rect 19810 3170 20390 3190
rect 19810 30 19830 3170
rect 20370 30 20390 3170
rect 19810 0 20390 30
rect 21010 3170 21590 3230
rect 21010 30 21030 3170
rect 21570 30 21590 3170
rect 21010 10 21590 30
rect 22210 3190 22790 3230
rect 22210 3170 23390 3190
rect 22210 30 22230 3170
rect 22770 30 22830 3170
rect 23370 30 23390 3170
rect 22210 10 23390 30
<< end >>
