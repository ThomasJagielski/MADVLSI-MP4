* SPICE3 file created from /home/madvlsi/Documents/MADVLSI-MP4/layout/ibias_vg.ext - technology: sky130A


* Top level circuit /home/madvlsi/Documents/MADVLSI-MP4/layout/ibias_vg

X0 a_15200_n14630# Vbn Vbp GND sky130_fd_pr__nfet_01v8 ad=1.28e+14p pd=8e+07u as=1.28e+14p ps=8e+07u w=1.6e+07u l=4e+06u
X1 Vr a_1600_n14660# a_1600_n14660# GND sky130_fd_pr__nfet_01v8 ad=3.84e+14p pd=2.4e+08u as=2.56e+14p ps=1.6e+08u w=1.6e+07u l=4e+06u
X2 net10 Vg VDD GND sky130_fd_pr__nfet_01v8 ad=1.28e+14p pd=8e+07u as=8.1987e+14p ps=6.061e+08u w=1.6e+07u l=4e+06u
X3 GND Vbn a_26400_n14630# GND sky130_fd_pr__nfet_01v8 ad=1.536e+15p pd=9.6e+08u as=1.28e+14p ps=8e+07u w=1.6e+07u l=4e+06u
X4 a_4000_n4790# Vbp VDD VDD sky130_fd_pr__pfet_01v8 ad=1.28e+14p pd=8e+07u as=1.28e+15p ps=8e+08u w=1.6e+07u l=4e+06u
X5 a_24800_n14630# GND GND GND sky130_fd_pr__nfet_01v8 ad=1.28e+14p pd=8e+07u as=0p ps=0u w=1.6e+07u l=4e+06u
X6 Vr GND GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X7 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X8 VDD Vg net13 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.28e+14p ps=8e+07u w=1.6e+07u l=4e+06u
X9 a_8800_n4790# Vdp Vdp VDD sky130_fd_pr__pfet_01v8 ad=1.28e+14p pd=8e+07u as=1.28e+14p ps=8e+07u w=1.6e+07u l=4e+06u
X10 GND GND GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X11 a_29600_n14630# net9 GND GND sky130_fd_pr__nfet_01v8 ad=1.28e+14p pd=8e+07u as=0p ps=0u w=1.6e+07u l=4e+06u
X12 a_29600_n14630# net9 GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X13 a_1600_n14660# a_1600_n14660# Vr GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X14 GND GND VDD GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X15 VDD Vdp a_8800_n4790# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X16 Vg a_24800_n14630# a_29600_n4790# VDD sky130_fd_pr__pfet_01v8 ad=1.28e+14p pd=8e+07u as=1.28e+14p ps=8e+07u w=1.6e+07u l=4e+06u
X17 Vdp a_1600_n14660# a_10400_n14630# GND sky130_fd_pr__nfet_01v8 ad=1.28e+14p pd=8e+07u as=1.28e+14p ps=8e+07u w=1.6e+07u l=4e+06u
X18 net11 Vg VDD GND sky130_fd_pr__nfet_01v8 ad=1.28e+14p pd=8e+07u as=0p ps=0u w=1.6e+07u l=4e+06u
X19 net9 Vg net11 GND sky130_fd_pr__nfet_01v8 ad=2.56e+14p pd=1.6e+08u as=0p ps=0u w=1.6e+07u l=4e+06u
X20 VDD Vbp a_16800_n4790# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.28e+14p ps=8e+07u w=1.6e+07u l=4e+06u
X21 Vbp GND Vdp GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X22 GND Vbn a_40000_n14630# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.28e+14p ps=8e+07u w=1.6e+07u l=4e+06u
X23 a_18400_n14630# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=1.28e+14p pd=8e+07u as=0p ps=0u w=1.6e+07u l=4e+06u
X24 Vbn VDD Vbp VDD sky130_fd_pr__pfet_01v8 ad=1.28e+14p pd=8e+07u as=1.28e+14p ps=8e+07u w=1.6e+07u l=4e+06u
X25 GND Vbn a_26400_n14630# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X26 a_1600_n14660# a_1600_n14660# Vr GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X27 a_12000_n4790# Vdp VDD VDD sky130_fd_pr__pfet_01v8 ad=1.28e+14p pd=8e+07u as=0p ps=0u w=1.6e+07u l=4e+06u
X28 Vr a_1600_n14660# a_1600_n14660# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X29 a_1600_n14660# Vbp a_4000_n4790# VDD sky130_fd_pr__pfet_01v8 ad=1.28e+14p pd=8e+07u as=0p ps=0u w=1.6e+07u l=4e+06u
X30 VDD Vg net10 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X31 Vbn VDD Vbp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X32 GND GND Vbn GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.28e+14p ps=8e+07u w=1.6e+07u l=4e+06u
X33 GND GND Vg GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.28e+14p ps=8e+07u w=1.6e+07u l=4e+06u
X34 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X35 Vg net9 a_29600_n14630# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X36 a_4000_n4790# Vbp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X37 a_24800_n14630# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=1.28e+14p pd=8e+07u as=0p ps=0u w=1.6e+07u l=4e+06u
X38 Vbn Vbn a_18400_n14630# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X39 GND GND VDD GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X40 net9 Vg net13 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X41 GND GND Vr GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X42 a_1600_n14660# Vbp a_4000_n4790# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X43 GND Vbn a_15200_n14630# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X44 a_26400_n4790# a_24800_n14630# a_24800_n14630# VDD sky130_fd_pr__pfet_01v8 ad=1.28e+14p pd=8e+07u as=0p ps=0u w=1.6e+07u l=4e+06u
X45 VDD a_24800_n14630# a_26400_n4790# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X46 a_24800_n14630# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X47 a_10400_n14630# a_1600_n14660# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X48 GND GND GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X49 VDD GND GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X50 VDD GND GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X51 Vr a_1600_n14660# a_1600_n14660# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X52 net9 Vbn a_40000_n14630# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X53 Vbp Vdp a_12000_n4790# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X54 a_15200_n14630# Vbn Vbp GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X55 net9 Vg net10 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X56 Vbn Vbn a_18400_n14630# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X57 a_24800_n14630# GND GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X58 Vr a_1600_n14660# a_1600_n14660# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X59 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X60 a_16800_n4790# Vbp Vbn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X61 Vbp GND Vdp GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X62 a_29600_n4790# a_24800_n14630# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X63 Vg a_24800_n14630# a_29600_n4790# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X64 VDD GND GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X65 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X66 a_26400_n14630# Vbn a_24800_n14630# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X67 a_1600_n14660# a_1600_n14660# Vr GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X68 VDD Vg net11 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X69 a_26400_n4790# a_24800_n14630# a_24800_n14630# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X70 GND GND Vg GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X71 VDD Vbp a_16800_n4790# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X72 net13 Vg net9 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X73 a_10400_n14630# a_1600_n14660# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X74 Vdp VDD a_1600_n14660# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X75 a_8800_n4790# Vdp Vdp VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X76 VDD a_24800_n14630# a_26400_n4790# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X77 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X78 Vdp a_1600_n14660# a_10400_n14630# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X79 Vr GND GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X80 net13 Vg VDD GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X81 a_29600_n4790# a_24800_n14630# VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X82 a_40000_n14630# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X83 GND GND Vr GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X84 a_40000_n14630# Vbn net9 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X85 a_12000_n4790# Vdp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X86 VDD VDD Vg VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X87 a_26400_n14630# Vbn a_24800_n14630# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X88 a_1600_n14660# a_1600_n14660# Vr GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X89 GND GND Vbn GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X90 GND GND VDD GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X91 GND Vbn a_15200_n14630# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X92 net10 Vg net9 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X93 Vbp Vdp a_12000_n4790# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X94 Vg net9 a_29600_n14630# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X95 net11 Vg net9 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X96 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X97 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X98 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X99 a_16800_n4790# Vbp Vbn VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X100 VDD Vdp a_8800_n4790# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X101 a_18400_n14630# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X102 VDD VDD Vg VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
X103 Vdp VDD a_1600_n14660# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.6e+07u l=4e+06u
.end

