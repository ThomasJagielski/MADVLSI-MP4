magic
tech sky130A
timestamp 1616796040
<< nwell >>
rect -190 -20 2810 170
<< pmos >>
rect 30 0 130 150
rect 230 0 330 150
rect 560 0 660 150
rect 760 0 860 150
rect 960 0 1060 150
rect 1160 0 1260 150
rect 1360 0 1460 150
rect 1560 0 1660 150
rect 1760 0 1860 150
rect 1960 0 2060 150
rect 2290 0 2390 150
rect 2490 0 2590 150
<< pdiff >>
rect -70 130 30 150
rect -70 20 -50 130
rect 10 20 30 130
rect -70 0 30 20
rect 130 130 230 150
rect 130 20 150 130
rect 210 20 230 130
rect 130 0 230 20
rect 330 130 430 150
rect 330 20 350 130
rect 410 20 430 130
rect 330 0 430 20
rect 460 130 560 150
rect 460 20 480 130
rect 540 20 560 130
rect 460 0 560 20
rect 660 130 760 150
rect 660 20 680 130
rect 740 20 760 130
rect 660 0 760 20
rect 860 130 960 150
rect 860 20 880 130
rect 940 20 960 130
rect 860 0 960 20
rect 1060 130 1160 150
rect 1060 20 1080 130
rect 1140 20 1160 130
rect 1060 0 1160 20
rect 1260 130 1360 150
rect 1260 20 1280 130
rect 1340 20 1360 130
rect 1260 0 1360 20
rect 1460 130 1560 150
rect 1460 20 1480 130
rect 1540 20 1560 130
rect 1460 0 1560 20
rect 1660 130 1760 150
rect 1660 20 1680 130
rect 1740 20 1760 130
rect 1660 0 1760 20
rect 1860 130 1960 150
rect 1860 20 1880 130
rect 1940 20 1960 130
rect 1860 0 1960 20
rect 2060 130 2160 150
rect 2060 20 2080 130
rect 2140 20 2160 130
rect 2060 0 2160 20
rect 2190 130 2290 150
rect 2190 20 2210 130
rect 2270 20 2290 130
rect 2190 0 2290 20
rect 2390 130 2490 150
rect 2390 20 2410 130
rect 2470 20 2490 130
rect 2390 0 2490 20
rect 2590 130 2690 150
rect 2590 20 2610 130
rect 2670 20 2690 130
rect 2590 0 2690 20
<< pdiffc >>
rect -50 20 10 130
rect 150 20 210 130
rect 350 20 410 130
rect 480 20 540 130
rect 680 20 740 130
rect 880 20 940 130
rect 1080 20 1140 130
rect 1280 20 1340 130
rect 1480 20 1540 130
rect 1680 20 1740 130
rect 1880 20 1940 130
rect 2080 20 2140 130
rect 2210 20 2270 130
rect 2410 20 2470 130
rect 2610 20 2670 130
<< nsubdiff >>
rect -170 130 -70 150
rect -170 20 -150 130
rect -90 20 -70 130
rect -170 0 -70 20
rect 2690 130 2790 150
rect 2690 20 2710 130
rect 2770 20 2790 130
rect 2690 0 2790 20
<< nsubdiffcont >>
rect -150 20 -90 130
rect 2710 20 2770 130
<< poly >>
rect 30 150 130 165
rect 230 150 330 165
rect 560 150 660 165
rect 760 150 860 165
rect 960 150 1060 165
rect 1160 150 1260 165
rect 1360 150 1460 165
rect 1560 150 1660 165
rect 1760 150 1860 165
rect 1960 150 2060 165
rect 2290 150 2390 165
rect 2490 150 2590 165
rect 30 -15 130 0
rect 230 -15 330 0
rect 560 -15 660 0
rect 760 -15 860 0
rect 960 -15 1060 0
rect 1160 -15 1260 0
rect 1360 -15 1460 0
rect 1560 -15 1660 0
rect 1760 -15 1860 0
rect 1960 -15 2060 0
rect 2290 -15 2390 0
rect 2490 -15 2590 0
rect 230 -25 660 -15
rect 230 -30 500 -25
rect 490 -45 500 -30
rect 520 -30 660 -25
rect 1960 -25 2390 -15
rect 1960 -30 2100 -25
rect 520 -45 530 -30
rect 490 -55 530 -45
rect 2090 -45 2100 -30
rect 2120 -30 2390 -25
rect 2120 -45 2130 -30
rect 2090 -55 2130 -45
<< polycont >>
rect 500 -45 520 -25
rect 2100 -45 2120 -25
<< locali >>
rect -160 130 20 140
rect -160 20 -150 130
rect -90 20 -50 130
rect 10 20 20 130
rect -160 10 20 20
rect 140 130 220 140
rect 140 20 150 130
rect 210 20 220 130
rect 140 10 220 20
rect 340 130 420 140
rect 340 20 350 130
rect 410 20 420 130
rect 340 10 420 20
rect 470 130 550 140
rect 470 20 480 130
rect 540 20 550 130
rect 470 10 550 20
rect 670 130 750 140
rect 670 20 680 130
rect 740 20 750 130
rect 670 10 750 20
rect 870 130 950 140
rect 870 20 880 130
rect 940 20 950 130
rect 870 10 950 20
rect 1070 130 1150 140
rect 1070 20 1080 130
rect 1140 20 1150 130
rect 1070 10 1150 20
rect 1270 130 1350 140
rect 1270 20 1280 130
rect 1340 20 1350 130
rect 1270 10 1350 20
rect 1470 130 1550 140
rect 1470 20 1480 130
rect 1540 20 1550 130
rect 1470 10 1550 20
rect 1670 130 1750 140
rect 1670 20 1680 130
rect 1740 20 1750 130
rect 1670 10 1750 20
rect 1870 130 1950 140
rect 1870 20 1880 130
rect 1940 20 1950 130
rect 1870 10 1950 20
rect 2070 130 2150 140
rect 2070 20 2080 130
rect 2140 20 2150 130
rect 2070 10 2150 20
rect 2200 130 2280 140
rect 2200 20 2210 130
rect 2270 20 2280 130
rect 2200 10 2280 20
rect 2400 130 2480 140
rect 2400 20 2410 130
rect 2470 20 2480 130
rect 2400 10 2480 20
rect 2600 130 2780 140
rect 2600 20 2610 130
rect 2670 20 2710 130
rect 2770 20 2780 130
rect 2600 10 2780 20
rect 490 -25 530 10
rect 490 -45 500 -25
rect 520 -45 530 -25
rect 490 -55 530 -45
rect 2090 -25 2130 10
rect 2090 -45 2100 -25
rect 2120 -45 2130 -25
rect 2090 -55 2130 -45
<< end >>
