magic
tech sky130A
timestamp 1617562696
<< nwell >>
rect 9225 160 9615 220
<< nmos >>
rect 5630 -7425 6030 -7420
rect 6430 -7425 6830 -7420
rect 8030 -7425 8430 -7420
rect 8830 -7425 9230 -7420
rect 10430 -7425 10830 -7420
rect 11230 -7425 11630 -7420
<< poly >>
rect 9225 205 9615 215
rect 9225 185 9235 205
rect 9605 185 9615 205
rect 9225 25 9615 185
rect 9225 5 9235 25
rect 9605 5 9615 25
rect 9225 -5 9615 5
rect 5630 -7460 6030 -7425
rect 5630 -7480 5640 -7460
rect 6020 -7480 6030 -7460
rect 5630 -7490 6030 -7480
rect 6430 -7460 6830 -7425
rect 6430 -7480 6440 -7460
rect 6820 -7480 6830 -7460
rect 6430 -7490 6830 -7480
rect 8030 -7460 8430 -7425
rect 8030 -7480 8040 -7460
rect 8420 -7480 8430 -7460
rect 8030 -7490 8430 -7480
rect 8830 -7460 9230 -7425
rect 8830 -7480 8840 -7460
rect 9220 -7480 9230 -7460
rect 8830 -7490 9230 -7480
rect 10430 -7460 10830 -7425
rect 10430 -7480 10440 -7460
rect 10820 -7480 10830 -7460
rect 10430 -7490 10830 -7480
rect 11230 -7460 11630 -7425
rect 11230 -7480 11240 -7460
rect 11620 -7480 11630 -7460
rect 11230 -7490 11630 -7480
<< polycont >>
rect 9235 185 9605 205
rect 9235 5 9605 25
rect 5640 -7480 6020 -7460
rect 6440 -7480 6820 -7460
rect 8040 -7480 8420 -7460
rect 8840 -7480 9220 -7460
rect 10440 -7480 10820 -7460
rect 11240 -7480 11620 -7460
<< locali >>
rect -675 330 -25 370
rect -65 140 -25 330
rect 9225 205 9615 280
rect 9225 185 9235 205
rect 9605 185 9615 205
rect 9225 175 9615 185
rect -65 120 0 140
rect 11645 100 12015 275
rect 11645 60 13625 100
rect 9225 25 12025 35
rect 9225 5 9235 25
rect 9605 5 12025 25
rect 9225 -5 12025 5
rect 11635 -1830 12025 -5
rect 13235 -1645 13625 60
rect -11280 -5440 -11260 -5435
rect -12900 -5735 -12860 -5475
rect -11300 -5735 -11260 -5440
rect -10500 -5735 -10460 -5435
rect -8900 -5735 -8860 -5460
rect -8100 -5735 -8060 -5470
rect -6500 -5735 -6460 -5470
rect -5700 -5735 -5660 -5470
rect 5630 -7460 6030 -7450
rect 5630 -7480 5640 -7460
rect 6020 -7480 6030 -7460
rect 5630 -7490 6030 -7480
rect 6430 -7460 6830 -7450
rect 6430 -7480 6440 -7460
rect 6820 -7480 6830 -7460
rect 6430 -7490 6830 -7480
rect 8030 -7460 8430 -7450
rect 8030 -7480 8040 -7460
rect 8420 -7480 8430 -7460
rect 8030 -7490 8430 -7480
rect 8830 -7460 9230 -7450
rect 8830 -7480 8840 -7460
rect 9220 -7480 9230 -7460
rect 8830 -7490 9230 -7480
rect 10430 -7460 10830 -7450
rect 10430 -7480 10440 -7460
rect 10820 -7480 10830 -7460
rect 10430 -7490 10830 -7480
rect 11230 -7460 11630 -7450
rect 11230 -7480 11240 -7460
rect 11620 -7480 11630 -7460
rect 11230 -7490 11630 -7480
<< viali >>
rect 4040 -7480 4420 -7460
rect 5640 -7480 6020 -7460
rect 6440 -7480 6820 -7460
rect 8040 -7480 8420 -7460
rect 8840 -7480 9220 -7460
rect 10440 -7480 10820 -7460
rect 11240 -7480 11620 -7460
<< metal1 >>
rect 4030 -7460 4430 -7420
rect 4030 -7480 4040 -7460
rect 4420 -7480 4430 -7460
rect 4030 -7490 4430 -7480
rect 5630 -7460 6030 -7420
rect 5630 -7480 5640 -7460
rect 6020 -7480 6030 -7460
rect 5630 -7490 6030 -7480
rect 6430 -7460 6830 -7420
rect 6430 -7480 6440 -7460
rect 6820 -7480 6830 -7460
rect 6430 -7490 6830 -7480
rect 8030 -7460 8430 -7420
rect 8030 -7480 8040 -7460
rect 8420 -7480 8430 -7460
rect 8030 -7490 8430 -7480
rect 8830 -7460 9230 -7420
rect 8830 -7480 8840 -7460
rect 9220 -7480 9230 -7460
rect 8830 -7490 9230 -7480
rect 10430 -7460 10830 -7420
rect 10430 -7480 10440 -7460
rect 10820 -7480 10830 -7460
rect 10430 -7490 10830 -7480
rect 11230 -7460 11630 -7420
rect 11230 -7480 11240 -7460
rect 11620 -7480 11630 -7460
rect 11230 -7490 11630 -7480
use mux2  mux2_6
timestamp 1616853209
transform 1 0 -5985 0 1 -6175
box 0 -60 415 505
use mux2  mux2_0
timestamp 1616853209
transform 1 0 -13185 0 1 -6175
box 0 -60 415 505
use dac_ladder  dac_ladder_1
timestamp 1617561611
transform 1 0 -12375 0 1 -1410
box -4700 -4135 11700 3405
use mux2  mux2_1
timestamp 1616853209
transform 1 0 -11585 0 1 -6175
box 0 -60 415 505
use mux2  mux2_2
timestamp 1616853209
transform 1 0 -10785 0 1 -6175
box 0 -60 415 505
use mux2  mux2_3
timestamp 1616853209
transform 1 0 -9185 0 1 -6175
box 0 -60 415 505
use mux2  mux2_4
timestamp 1616853209
transform 1 0 -8385 0 1 -6175
box 0 -60 415 505
use mux2  mux2_5
timestamp 1616853209
transform 1 0 -6785 0 1 -6175
box 0 -60 415 505
use low-voltage_super-wilson  low-voltage_super-wilson_0
timestamp 1617552636
transform 1 0 615 0 1 275
box -615 -275 15825 1785
use dac_ladder  dac_ladder_0
timestamp 1617561611
transform 1 0 4730 0 1 -3425
box -4700 -4135 11700 3405
use ibias_vg  ibias_vg_0
timestamp 1617552423
transform 1 0 -16090 0 1 10945
box -820 -8300 24030 2600
<< labels >>
rlabel poly 5885 -7490 5885 -7490 5 b0
rlabel poly 6685 -7490 6685 -7490 5 b0
rlabel poly 8285 -7490 8285 -7490 5 b0
rlabel poly 9085 -7490 9085 -7490 5 b0
rlabel poly 10685 -7490 10685 -7490 5 b0
rlabel poly 11485 -7490 11485 -7490 5 b0
<< end >>
