magic
tech sky130A
timestamp 1616836363
<< nwell >>
rect -190 -20 250 170
rect -190 -520 250 -330
<< pwell >>
rect -190 -1020 250 -830
<< nmos >>
rect 30 -1000 130 -850
<< pmos >>
rect 30 0 130 150
rect 30 -500 130 -350
<< ndiff >>
rect -70 -870 30 -850
rect -70 -980 -50 -870
rect 10 -980 30 -870
rect -70 -1000 30 -980
rect 130 -870 230 -850
rect 130 -980 150 -870
rect 210 -980 230 -870
rect 130 -1000 230 -980
<< pdiff >>
rect -70 130 30 150
rect -70 20 -50 130
rect 10 20 30 130
rect -70 0 30 20
rect 130 130 230 150
rect 130 20 150 130
rect 210 20 230 130
rect 130 0 230 20
rect -70 -370 30 -350
rect -70 -480 -50 -370
rect 10 -480 30 -370
rect -70 -500 30 -480
rect 130 -370 230 -350
rect 130 -480 150 -370
rect 210 -480 230 -370
rect 130 -500 230 -480
<< ndiffc >>
rect -50 -980 10 -870
rect 150 -980 210 -870
<< pdiffc >>
rect -50 20 10 130
rect 150 20 210 130
rect -50 -480 10 -370
rect 150 -480 210 -370
<< psubdiff >>
rect -170 -870 -70 -850
rect -170 -980 -150 -870
rect -90 -980 -70 -870
rect -170 -1000 -70 -980
<< nsubdiff >>
rect -170 130 -70 150
rect -170 20 -150 130
rect -90 20 -70 130
rect -170 0 -70 20
rect -170 -370 -70 -350
rect -170 -480 -150 -370
rect -90 -480 -70 -370
rect -170 -500 -70 -480
<< psubdiffcont >>
rect -150 -980 -90 -870
<< nsubdiffcont >>
rect -150 20 -90 130
rect -150 -480 -90 -370
<< poly >>
rect 30 150 130 165
rect 30 -15 130 0
rect 30 -350 130 -335
rect 30 -515 130 -500
rect 30 -850 130 -835
rect 30 -1015 130 -1000
<< locali >>
rect -160 130 20 140
rect -160 20 -150 130
rect -90 20 -50 130
rect 10 20 20 130
rect -160 10 20 20
rect 140 130 220 140
rect 140 20 150 130
rect 210 20 220 130
rect 140 10 220 20
rect -160 -370 20 -360
rect -160 -480 -150 -370
rect -90 -480 -50 -370
rect 10 -480 20 -370
rect -160 -490 20 -480
rect 140 -370 220 -360
rect 140 -480 150 -370
rect 210 -480 220 -370
rect 140 -490 220 -480
rect -160 -870 20 -860
rect -160 -980 -150 -870
rect -90 -980 -50 -870
rect 10 -980 20 -870
rect -160 -990 20 -980
rect 140 -870 220 -860
rect 140 -980 150 -870
rect 210 -980 220 -870
rect 140 -990 220 -980
<< end >>
