magic
tech sky130A
timestamp 1616837863
<< error_p >>
rect 1430 0 1530 150
<< nwell >>
rect -190 -20 3150 170
<< pmos >>
rect 30 0 130 150
rect 230 0 330 150
rect 430 0 530 150
rect 630 0 730 150
rect 755 0 855 150
rect 880 0 980 150
rect 1005 0 1105 150
rect 1130 0 1230 150
rect 1330 0 1430 150
rect 1530 0 1630 150
rect 1730 0 1830 150
rect 1855 0 1955 150
rect 1980 0 2080 150
rect 2105 0 2205 150
rect 2230 0 2330 150
rect 2430 0 2530 150
rect 2630 0 2730 150
rect 2830 0 2930 150
<< pdiff >>
rect -70 130 30 150
rect -70 20 -50 130
rect 10 20 30 130
rect -70 0 30 20
rect 130 130 230 150
rect 130 20 150 130
rect 210 20 230 130
rect 130 0 230 20
rect 330 130 430 150
rect 330 20 350 130
rect 410 20 430 130
rect 330 0 430 20
rect 530 130 630 150
rect 530 20 550 130
rect 610 20 630 130
rect 530 0 630 20
rect 730 0 755 150
rect 855 0 880 150
rect 980 0 1005 150
rect 1105 0 1130 150
rect 1230 130 1330 150
rect 1230 20 1250 130
rect 1310 20 1330 130
rect 1230 0 1330 20
rect 1430 130 1530 150
rect 1430 20 1450 130
rect 1510 20 1530 130
rect 1430 0 1530 20
rect 1630 130 1730 150
rect 1630 20 1650 130
rect 1710 20 1730 130
rect 1630 0 1730 20
rect 1830 0 1855 150
rect 1955 0 1980 150
rect 2080 0 2105 150
rect 2205 0 2230 150
rect 2330 130 2430 150
rect 2330 20 2350 130
rect 2410 20 2430 130
rect 2330 0 2430 20
rect 2530 130 2630 150
rect 2530 20 2550 130
rect 2610 20 2630 130
rect 2530 0 2630 20
rect 2730 130 2830 150
rect 2730 20 2750 130
rect 2810 20 2830 130
rect 2730 0 2830 20
rect 2930 130 3030 150
rect 2930 20 2950 130
rect 3010 20 3030 130
rect 2930 0 3030 20
<< pdiffc >>
rect -50 20 10 130
rect 150 20 210 130
rect 350 20 410 130
rect 550 20 610 130
rect 1250 20 1310 130
rect 1450 20 1510 130
rect 1650 20 1710 130
rect 2350 20 2410 130
rect 2550 20 2610 130
rect 2750 20 2810 130
rect 2950 20 3010 130
<< nsubdiff >>
rect -170 130 -70 150
rect -170 20 -150 130
rect -90 20 -70 130
rect -170 0 -70 20
rect 3030 130 3130 150
rect 3030 20 3050 130
rect 3110 20 3130 130
rect 3030 0 3130 20
<< nsubdiffcont >>
rect -150 20 -90 130
rect 3050 20 3110 130
<< poly >>
rect 30 150 130 165
rect 230 150 330 165
rect 430 150 530 165
rect 630 150 730 165
rect 755 150 855 165
rect 880 150 980 165
rect 1005 150 1105 165
rect 1130 150 1230 165
rect 1330 150 1430 165
rect 1530 150 1630 165
rect 1730 150 1830 165
rect 1855 150 1955 165
rect 1980 150 2080 165
rect 2105 150 2205 165
rect 2230 150 2330 165
rect 2430 150 2530 165
rect 2630 150 2730 165
rect 2830 150 2930 165
rect 30 -15 130 0
rect 230 -15 330 0
rect 430 -15 530 0
rect 630 -15 730 0
rect 755 -15 855 0
rect 880 -15 980 0
rect 1005 -15 1105 0
rect 1130 -15 1230 0
rect 1330 -15 1430 0
rect 1530 -15 1630 0
rect 1730 -15 1830 0
rect 1855 -15 1955 0
rect 1980 -15 2080 0
rect 2105 -15 2205 0
rect 2230 -15 2330 0
rect 2430 -15 2530 0
rect 2630 -15 2730 0
rect 2830 -15 2930 0
<< locali >>
rect -160 130 20 140
rect -160 20 -150 130
rect -90 20 -50 130
rect 10 20 20 130
rect -160 10 20 20
rect 140 130 220 140
rect 140 20 150 130
rect 210 20 220 130
rect 140 10 220 20
rect 340 130 420 140
rect 340 20 350 130
rect 410 20 420 130
rect 340 10 420 20
rect 540 130 620 140
rect 540 20 550 130
rect 610 20 620 130
rect 540 10 620 20
rect 1240 130 1320 140
rect 1240 20 1250 130
rect 1310 20 1320 130
rect 1240 10 1320 20
rect 1440 130 1520 140
rect 1440 20 1450 130
rect 1510 20 1520 130
rect 1440 10 1520 20
rect 1640 130 1720 140
rect 1640 20 1650 130
rect 1710 20 1720 130
rect 1640 10 1720 20
rect 2340 130 2420 140
rect 2340 20 2350 130
rect 2410 20 2420 130
rect 2340 10 2420 20
rect 2540 130 2620 140
rect 2540 20 2550 130
rect 2610 20 2620 130
rect 2540 10 2620 20
rect 2740 130 2820 140
rect 2740 20 2750 130
rect 2810 20 2820 130
rect 2740 10 2820 20
rect 2940 130 3120 140
rect 2940 20 2950 130
rect 3010 20 3050 130
rect 3110 20 3120 130
rect 2940 10 3120 20
<< end >>
