magic
tech sky130A
timestamp 1616853209
<< nwell >>
rect 135 230 415 470
<< nmos >>
rect 265 15 280 115
rect 330 15 345 115
<< pmos >>
rect 265 345 280 445
rect 330 345 345 445
<< ndiff >>
rect 215 100 265 115
rect 215 30 230 100
rect 250 30 265 100
rect 215 15 265 30
rect 280 100 330 115
rect 280 30 295 100
rect 315 30 330 100
rect 280 15 330 30
rect 345 100 395 115
rect 345 30 360 100
rect 380 30 395 100
rect 345 15 395 30
<< pdiff >>
rect 215 430 265 445
rect 215 360 230 430
rect 250 360 265 430
rect 215 345 265 360
rect 280 430 330 445
rect 280 360 295 430
rect 315 360 330 430
rect 280 345 330 360
rect 345 430 395 445
rect 345 360 360 430
rect 380 360 395 430
rect 345 345 395 360
<< ndiffc >>
rect 230 30 250 100
rect 295 30 315 100
rect 360 30 380 100
<< pdiffc >>
rect 230 360 250 430
rect 295 360 315 430
rect 360 360 380 430
<< poly >>
rect 135 490 345 505
rect 265 445 280 460
rect 330 445 345 490
rect 265 230 280 345
rect 330 330 345 345
rect 160 220 345 230
rect 160 200 170 220
rect 190 215 345 220
rect 190 200 200 215
rect 160 190 200 200
rect 120 125 280 140
rect 265 115 280 125
rect 330 115 345 215
rect 265 0 280 15
rect 330 0 345 15
<< polycont >>
rect 170 200 190 220
<< locali >>
rect 0 485 15 505
rect 305 485 415 505
rect 305 440 325 485
rect 220 430 260 440
rect 220 360 230 430
rect 250 360 260 430
rect 220 350 260 360
rect 285 430 325 440
rect 285 360 295 430
rect 315 360 325 430
rect 285 350 325 360
rect 350 430 390 440
rect 350 360 360 430
rect 380 360 390 430
rect 350 350 390 360
rect 160 220 200 230
rect 160 200 170 220
rect 190 200 200 220
rect 160 190 200 200
rect 220 110 240 350
rect 285 110 305 350
rect 350 110 370 350
rect 220 100 260 110
rect 220 30 230 100
rect 250 30 260 100
rect 220 20 260 30
rect 285 100 325 110
rect 285 30 295 100
rect 315 30 325 100
rect 285 20 325 30
rect 350 100 390 110
rect 350 30 360 100
rect 380 30 390 100
rect 350 20 390 30
rect 220 0 240 20
rect 0 -20 240 0
rect 350 -40 370 20
rect 0 -60 370 -40
<< metal1 >>
rect 0 255 20 445
rect 205 255 415 445
rect 0 20 20 210
rect 205 20 415 210
use inverter  inverter_0
timestamp 1616851029
transform 1 0 120 0 1 -120
box -120 120 85 625
<< labels >>
rlabel locali 415 495 415 495 3 muxout
rlabel locali 0 -10 0 -10 7 A
rlabel locali 0 -50 0 -50 7 B
rlabel locali 0 495 0 495 7 S
rlabel metal1 0 350 0 350 7 VP
rlabel metal1 0 115 0 115 7 VN
<< end >>
