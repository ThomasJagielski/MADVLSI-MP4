magic
tech sky130A
timestamp 1617392463
<< error_p >>
rect 20000 5 20400 1605
rect 20800 5 21200 1605
rect 21600 5 22000 1605
rect 20000 -2395 20400 -795
rect 20800 -2395 21200 -795
rect 21600 -2395 22000 -795
rect 20000 -4915 20400 -3315
rect 20800 -4915 21200 -3315
rect 21600 -4915 22000 -3315
rect 20000 -7315 20400 -5715
rect 20800 -7315 21200 -5715
rect 21600 -7315 22000 -5715
<< nmos >>
rect 0 5 400 1605
rect 800 5 1200 1605
rect 1600 5 2000 1605
rect 2400 5 2800 1605
rect 3200 5 3600 1605
rect 4000 5 4400 1605
rect 4800 5 5200 1605
rect 5600 5 6000 1605
rect 6400 5 6800 1605
rect 7200 5 7600 1605
rect 8000 5 8400 1605
rect 8800 5 9200 1605
rect 9600 5 10000 1605
rect 10400 5 10800 1605
rect 12000 5 12400 1605
rect 12800 5 13200 1605
rect 13600 5 14000 1605
rect 14400 5 14800 1605
rect 15200 5 15600 1605
rect 16000 5 16400 1605
rect 18800 5 19200 1605
rect 19600 5 20000 1605
rect 20400 5 20800 1605
rect 21200 5 21600 1605
rect 22000 5 22400 1605
rect 22800 5 23200 1605
rect 0 -2395 400 -795
rect 800 -2395 1200 -795
rect 1600 -2395 2000 -795
rect 2400 -2395 2800 -795
rect 3200 -2395 3600 -795
rect 4000 -2395 4400 -795
rect 4800 -2395 5200 -795
rect 5600 -2395 6000 -795
rect 6400 -2395 6800 -795
rect 7200 -2395 7600 -795
rect 8000 -2395 8400 -795
rect 8800 -2395 9200 -795
rect 9600 -2395 10000 -795
rect 10400 -2395 10800 -795
rect 12000 -2395 12400 -795
rect 12800 -2395 13200 -795
rect 13600 -2395 14000 -795
rect 14400 -2395 14800 -795
rect 15200 -2395 15600 -795
rect 16000 -2395 16400 -795
rect 18800 -2395 19200 -795
rect 19600 -2395 20000 -795
rect 20400 -2395 20800 -795
rect 21200 -2395 21600 -795
rect 22000 -2395 22400 -795
rect 22800 -2395 23200 -795
rect 0 -4915 400 -3315
rect 800 -4915 1200 -3315
rect 1600 -4915 2000 -3315
rect 2400 -4915 2800 -3315
rect 3200 -4915 3600 -3315
rect 4000 -4915 4400 -3315
rect 4800 -4915 5200 -3315
rect 5600 -4915 6000 -3315
rect 6400 -4915 6800 -3315
rect 7200 -4915 7600 -3315
rect 8000 -4915 8400 -3315
rect 8800 -4915 9200 -3315
rect 9600 -4915 10000 -3315
rect 10400 -4915 10800 -3315
rect 12000 -4915 12400 -3315
rect 12800 -4915 13200 -3315
rect 13600 -4915 14000 -3315
rect 14400 -4915 14800 -3315
rect 15200 -4915 15600 -3315
rect 16000 -4915 16400 -3315
rect 18800 -4915 19200 -3315
rect 19600 -4915 20000 -3315
rect 20400 -4915 20800 -3315
rect 21200 -4915 21600 -3315
rect 22000 -4915 22400 -3315
rect 22800 -4915 23200 -3315
rect 0 -7315 400 -5715
rect 800 -7315 1200 -5715
rect 1600 -7315 2000 -5715
rect 2400 -7315 2800 -5715
rect 3200 -7315 3600 -5715
rect 4000 -7315 4400 -5715
rect 4800 -7315 5200 -5715
rect 5600 -7315 6000 -5715
rect 6400 -7315 6800 -5715
rect 7200 -7315 7600 -5715
rect 8000 -7315 8400 -5715
rect 8800 -7315 9200 -5715
rect 9600 -7315 10000 -5715
rect 10400 -7315 10800 -5715
rect 12000 -7315 12400 -5715
rect 12800 -7315 13200 -5715
rect 13600 -7315 14000 -5715
rect 14400 -7315 14800 -5715
rect 15200 -7315 15600 -5715
rect 16000 -7315 16400 -5715
rect 18800 -7315 19200 -5715
rect 19600 -7315 20000 -5715
rect 20400 -7315 20800 -5715
rect 21200 -7315 21600 -5715
rect 22000 -7315 22400 -5715
rect 22800 -7315 23200 -5715
<< ndiff >>
rect -400 1585 0 1605
rect -400 25 -380 1585
rect -20 25 0 1585
rect -400 5 0 25
rect 400 1585 800 1605
rect 400 25 420 1585
rect 780 25 800 1585
rect 400 5 800 25
rect 1200 1585 1600 1605
rect 1200 25 1220 1585
rect 1580 25 1600 1585
rect 1200 5 1600 25
rect 2000 1585 2400 1605
rect 2000 25 2020 1585
rect 2380 25 2400 1585
rect 2000 5 2400 25
rect 2800 1585 3200 1605
rect 2800 25 2820 1585
rect 3180 25 3200 1585
rect 2800 5 3200 25
rect 3600 1585 4000 1605
rect 3600 25 3620 1585
rect 3980 25 4000 1585
rect 3600 5 4000 25
rect 4400 1585 4800 1605
rect 4400 25 4420 1585
rect 4780 25 4800 1585
rect 4400 5 4800 25
rect 5200 1585 5600 1605
rect 5200 25 5220 1585
rect 5580 25 5600 1585
rect 5200 5 5600 25
rect 6000 1585 6400 1605
rect 6000 25 6020 1585
rect 6380 25 6400 1585
rect 6000 5 6400 25
rect 6800 1585 7200 1605
rect 6800 25 6820 1585
rect 7180 25 7200 1585
rect 6800 5 7200 25
rect 7600 1585 8000 1605
rect 7600 25 7620 1585
rect 7980 25 8000 1585
rect 7600 5 8000 25
rect 8400 1585 8800 1605
rect 8400 25 8420 1585
rect 8780 25 8800 1585
rect 8400 5 8800 25
rect 9200 1585 9600 1605
rect 9200 25 9220 1585
rect 9580 25 9600 1585
rect 9200 5 9600 25
rect 10000 1585 10400 1605
rect 10000 25 10020 1585
rect 10380 25 10400 1585
rect 10000 5 10400 25
rect 10800 1585 11200 1605
rect 11600 1585 12000 1605
rect 10800 25 10820 1585
rect 11180 25 11200 1585
rect 11600 25 11620 1585
rect 11980 25 12000 1585
rect 10800 5 11200 25
rect 11600 5 12000 25
rect 12400 1585 12800 1605
rect 12400 25 12420 1585
rect 12780 25 12800 1585
rect 12400 5 12800 25
rect 13200 1585 13600 1605
rect 13200 25 13220 1585
rect 13580 25 13600 1585
rect 13200 5 13600 25
rect 14000 1585 14400 1605
rect 14000 25 14020 1585
rect 14380 25 14400 1585
rect 14000 5 14400 25
rect 14800 1585 15200 1605
rect 14800 25 14820 1585
rect 15180 25 15200 1585
rect 14800 5 15200 25
rect 15600 1585 16000 1605
rect 15600 25 15620 1585
rect 15980 25 16000 1585
rect 15600 5 16000 25
rect 16400 1585 16800 1605
rect 16400 25 16420 1585
rect 16780 25 16800 1585
rect 16400 5 16800 25
rect 18400 1585 18800 1605
rect 18400 25 18420 1585
rect 18780 25 18800 1585
rect 18400 5 18800 25
rect 19200 1585 19600 1605
rect 19200 25 19220 1585
rect 19580 25 19600 1585
rect 19200 5 19600 25
rect 20000 1585 20400 1605
rect 20000 25 20020 1585
rect 20380 25 20400 1585
rect 20000 5 20400 25
rect 20800 1585 21200 1605
rect 20800 25 20820 1585
rect 21180 25 21200 1585
rect 20800 5 21200 25
rect 21600 1585 22000 1605
rect 21600 25 21620 1585
rect 21980 25 22000 1585
rect 21600 5 22000 25
rect 22400 1585 22800 1605
rect 22400 25 22420 1585
rect 22780 25 22800 1585
rect 22400 5 22800 25
rect 23200 1585 23600 1605
rect 23200 25 23220 1585
rect 23580 25 23600 1585
rect 23200 5 23600 25
rect -400 -815 0 -795
rect -400 -2375 -380 -815
rect -20 -2375 0 -815
rect -400 -2395 0 -2375
rect 400 -815 800 -795
rect 400 -2375 420 -815
rect 780 -2375 800 -815
rect 400 -2395 800 -2375
rect 1200 -815 1600 -795
rect 1200 -2375 1220 -815
rect 1580 -2375 1600 -815
rect 1200 -2395 1600 -2375
rect 2000 -815 2400 -795
rect 2000 -2375 2020 -815
rect 2380 -2375 2400 -815
rect 2000 -2395 2400 -2375
rect 2800 -815 3200 -795
rect 2800 -2375 2820 -815
rect 3180 -2375 3200 -815
rect 2800 -2395 3200 -2375
rect 3600 -815 4000 -795
rect 3600 -2375 3620 -815
rect 3980 -2375 4000 -815
rect 3600 -2395 4000 -2375
rect 4400 -815 4800 -795
rect 4400 -2375 4420 -815
rect 4780 -2375 4800 -815
rect 4400 -2395 4800 -2375
rect 5200 -815 5600 -795
rect 5200 -2375 5220 -815
rect 5580 -2375 5600 -815
rect 5200 -2395 5600 -2375
rect 6000 -815 6400 -795
rect 6000 -2375 6020 -815
rect 6380 -2375 6400 -815
rect 6000 -2395 6400 -2375
rect 6800 -815 7200 -795
rect 6800 -2375 6820 -815
rect 7180 -2375 7200 -815
rect 6800 -2395 7200 -2375
rect 7600 -815 8000 -795
rect 7600 -2375 7620 -815
rect 7980 -2375 8000 -815
rect 7600 -2395 8000 -2375
rect 8400 -815 8800 -795
rect 8400 -2375 8420 -815
rect 8780 -2375 8800 -815
rect 8400 -2395 8800 -2375
rect 9200 -815 9600 -795
rect 9200 -2375 9220 -815
rect 9580 -2375 9600 -815
rect 9200 -2395 9600 -2375
rect 10000 -815 10400 -795
rect 10000 -2375 10020 -815
rect 10380 -2375 10400 -815
rect 10000 -2395 10400 -2375
rect 10800 -815 11200 -795
rect 11600 -815 12000 -795
rect 10800 -2375 10820 -815
rect 11180 -2375 11200 -815
rect 11600 -2375 11620 -815
rect 11980 -2375 12000 -815
rect 10800 -2395 11200 -2375
rect 11600 -2395 12000 -2375
rect 12400 -815 12800 -795
rect 12400 -2375 12420 -815
rect 12780 -2375 12800 -815
rect 12400 -2395 12800 -2375
rect 13200 -815 13600 -795
rect 13200 -2375 13220 -815
rect 13580 -2375 13600 -815
rect 13200 -2395 13600 -2375
rect 14000 -815 14400 -795
rect 14000 -2375 14020 -815
rect 14380 -2375 14400 -815
rect 14000 -2395 14400 -2375
rect 14800 -815 15200 -795
rect 14800 -2375 14820 -815
rect 15180 -2375 15200 -815
rect 14800 -2395 15200 -2375
rect 15600 -815 16000 -795
rect 15600 -2375 15620 -815
rect 15980 -2375 16000 -815
rect 15600 -2395 16000 -2375
rect 16400 -815 16800 -795
rect 16400 -2375 16420 -815
rect 16780 -2375 16800 -815
rect 16400 -2395 16800 -2375
rect 18400 -815 18800 -795
rect 18400 -2375 18420 -815
rect 18780 -2375 18800 -815
rect 18400 -2395 18800 -2375
rect 19200 -815 19600 -795
rect 19200 -2375 19220 -815
rect 19580 -2375 19600 -815
rect 19200 -2395 19600 -2375
rect 20000 -815 20400 -795
rect 20000 -2375 20020 -815
rect 20380 -2375 20400 -815
rect 20000 -2395 20400 -2375
rect 20800 -815 21200 -795
rect 20800 -2375 20820 -815
rect 21180 -2375 21200 -815
rect 20800 -2395 21200 -2375
rect 21600 -815 22000 -795
rect 21600 -2375 21620 -815
rect 21980 -2375 22000 -815
rect 21600 -2395 22000 -2375
rect 22400 -815 22800 -795
rect 22400 -2375 22420 -815
rect 22780 -2375 22800 -815
rect 22400 -2395 22800 -2375
rect 23200 -815 23600 -795
rect 23200 -2375 23220 -815
rect 23580 -2375 23600 -815
rect 23200 -2395 23600 -2375
rect -400 -3335 0 -3315
rect -400 -4895 -380 -3335
rect -20 -4895 0 -3335
rect -400 -4915 0 -4895
rect 400 -3335 800 -3315
rect 400 -4895 420 -3335
rect 780 -4895 800 -3335
rect 400 -4915 800 -4895
rect 1200 -3335 1600 -3315
rect 1200 -4895 1220 -3335
rect 1580 -4895 1600 -3335
rect 1200 -4915 1600 -4895
rect 2000 -3335 2400 -3315
rect 2000 -4895 2020 -3335
rect 2380 -4895 2400 -3335
rect 2000 -4915 2400 -4895
rect 2800 -3335 3200 -3315
rect 2800 -4895 2820 -3335
rect 3180 -4895 3200 -3335
rect 2800 -4915 3200 -4895
rect 3600 -3335 4000 -3315
rect 3600 -4895 3620 -3335
rect 3980 -4895 4000 -3335
rect 3600 -4915 4000 -4895
rect 4400 -3335 4800 -3315
rect 4400 -4895 4420 -3335
rect 4780 -4895 4800 -3335
rect 4400 -4915 4800 -4895
rect 5200 -3335 5600 -3315
rect 5200 -4895 5220 -3335
rect 5580 -4895 5600 -3335
rect 5200 -4915 5600 -4895
rect 6000 -3335 6400 -3315
rect 6000 -4895 6020 -3335
rect 6380 -4895 6400 -3335
rect 6000 -4915 6400 -4895
rect 6800 -3335 7200 -3315
rect 6800 -4895 6820 -3335
rect 7180 -4895 7200 -3335
rect 6800 -4915 7200 -4895
rect 7600 -3335 8000 -3315
rect 7600 -4895 7620 -3335
rect 7980 -4895 8000 -3335
rect 7600 -4915 8000 -4895
rect 8400 -3335 8800 -3315
rect 8400 -4895 8420 -3335
rect 8780 -4895 8800 -3335
rect 8400 -4915 8800 -4895
rect 9200 -3335 9600 -3315
rect 9200 -4895 9220 -3335
rect 9580 -4895 9600 -3335
rect 9200 -4915 9600 -4895
rect 10000 -3335 10400 -3315
rect 10000 -4895 10020 -3335
rect 10380 -4895 10400 -3335
rect 10000 -4915 10400 -4895
rect 10800 -3335 11200 -3315
rect 11600 -3335 12000 -3315
rect 10800 -4895 10820 -3335
rect 11180 -4895 11200 -3335
rect 11600 -4895 11620 -3335
rect 11980 -4895 12000 -3335
rect 10800 -4915 11200 -4895
rect 11600 -4915 12000 -4895
rect 12400 -3335 12800 -3315
rect 12400 -4895 12420 -3335
rect 12780 -4895 12800 -3335
rect 12400 -4915 12800 -4895
rect 13200 -3335 13600 -3315
rect 13200 -4895 13220 -3335
rect 13580 -4895 13600 -3335
rect 13200 -4915 13600 -4895
rect 14000 -3335 14400 -3315
rect 14000 -4895 14020 -3335
rect 14380 -4895 14400 -3335
rect 14000 -4915 14400 -4895
rect 14800 -3335 15200 -3315
rect 14800 -4895 14820 -3335
rect 15180 -4895 15200 -3335
rect 14800 -4915 15200 -4895
rect 15600 -3335 16000 -3315
rect 15600 -4895 15620 -3335
rect 15980 -4895 16000 -3335
rect 15600 -4915 16000 -4895
rect 16400 -3335 16800 -3315
rect 16400 -4895 16420 -3335
rect 16780 -4895 16800 -3335
rect 16400 -4915 16800 -4895
rect 18400 -3335 18800 -3315
rect 18400 -4895 18420 -3335
rect 18780 -4895 18800 -3335
rect 18400 -4915 18800 -4895
rect 19200 -3335 19600 -3315
rect 19200 -4895 19220 -3335
rect 19580 -4895 19600 -3335
rect 19200 -4915 19600 -4895
rect 20000 -3335 20400 -3315
rect 20000 -4895 20020 -3335
rect 20380 -4895 20400 -3335
rect 20000 -4915 20400 -4895
rect 20800 -3335 21200 -3315
rect 20800 -4895 20820 -3335
rect 21180 -4895 21200 -3335
rect 20800 -4915 21200 -4895
rect 21600 -3335 22000 -3315
rect 21600 -4895 21620 -3335
rect 21980 -4895 22000 -3335
rect 21600 -4915 22000 -4895
rect 22400 -3335 22800 -3315
rect 22400 -4895 22420 -3335
rect 22780 -4895 22800 -3335
rect 22400 -4915 22800 -4895
rect 23200 -3335 23600 -3315
rect 23200 -4895 23220 -3335
rect 23580 -4895 23600 -3335
rect 23200 -4915 23600 -4895
rect -400 -5735 0 -5715
rect -400 -7295 -380 -5735
rect -20 -7295 0 -5735
rect -400 -7315 0 -7295
rect 400 -5735 800 -5715
rect 400 -7295 420 -5735
rect 780 -7295 800 -5735
rect 400 -7315 800 -7295
rect 1200 -5735 1600 -5715
rect 1200 -7295 1220 -5735
rect 1580 -7295 1600 -5735
rect 1200 -7315 1600 -7295
rect 2000 -5735 2400 -5715
rect 2000 -7295 2020 -5735
rect 2380 -7295 2400 -5735
rect 2000 -7315 2400 -7295
rect 2800 -5735 3200 -5715
rect 2800 -7295 2820 -5735
rect 3180 -7295 3200 -5735
rect 2800 -7315 3200 -7295
rect 3600 -5735 4000 -5715
rect 3600 -7295 3620 -5735
rect 3980 -7295 4000 -5735
rect 3600 -7315 4000 -7295
rect 4400 -5735 4800 -5715
rect 4400 -7295 4420 -5735
rect 4780 -7295 4800 -5735
rect 4400 -7315 4800 -7295
rect 5200 -5735 5600 -5715
rect 5200 -7295 5220 -5735
rect 5580 -7295 5600 -5735
rect 5200 -7315 5600 -7295
rect 6000 -5735 6400 -5715
rect 6000 -7295 6020 -5735
rect 6380 -7295 6400 -5735
rect 6000 -7315 6400 -7295
rect 6800 -5735 7200 -5715
rect 6800 -7295 6820 -5735
rect 7180 -7295 7200 -5735
rect 6800 -7315 7200 -7295
rect 7600 -5735 8000 -5715
rect 7600 -7295 7620 -5735
rect 7980 -7295 8000 -5735
rect 7600 -7315 8000 -7295
rect 8400 -5735 8800 -5715
rect 8400 -7295 8420 -5735
rect 8780 -7295 8800 -5735
rect 8400 -7315 8800 -7295
rect 9200 -5735 9600 -5715
rect 9200 -7295 9220 -5735
rect 9580 -7295 9600 -5735
rect 9200 -7315 9600 -7295
rect 10000 -5735 10400 -5715
rect 10000 -7295 10020 -5735
rect 10380 -7295 10400 -5735
rect 10000 -7315 10400 -7295
rect 10800 -5735 11200 -5715
rect 11600 -5735 12000 -5715
rect 10800 -7295 10820 -5735
rect 11180 -7295 11200 -5735
rect 11600 -7295 11620 -5735
rect 11980 -7295 12000 -5735
rect 10800 -7315 11200 -7295
rect 11600 -7315 12000 -7295
rect 12400 -5735 12800 -5715
rect 12400 -7295 12420 -5735
rect 12780 -7295 12800 -5735
rect 12400 -7315 12800 -7295
rect 13200 -5735 13600 -5715
rect 13200 -7295 13220 -5735
rect 13580 -7295 13600 -5735
rect 13200 -7315 13600 -7295
rect 14000 -5735 14400 -5715
rect 14000 -7295 14015 -5735
rect 14380 -7295 14400 -5735
rect 14000 -7315 14400 -7295
rect 14800 -5735 15200 -5715
rect 14800 -7295 14820 -5735
rect 15180 -7295 15200 -5735
rect 14800 -7315 15200 -7295
rect 15600 -5735 16000 -5715
rect 15600 -7295 15620 -5735
rect 15980 -7295 16000 -5735
rect 15600 -7315 16000 -7295
rect 16400 -5735 16800 -5715
rect 16400 -7295 16420 -5735
rect 16780 -7295 16800 -5735
rect 16400 -7315 16800 -7295
rect 18400 -5735 18800 -5715
rect 18400 -7295 18420 -5735
rect 18780 -7295 18800 -5735
rect 18400 -7315 18800 -7295
rect 19200 -5735 19600 -5715
rect 19200 -7295 19220 -5735
rect 19580 -7295 19600 -5735
rect 19200 -7315 19600 -7295
rect 20000 -5735 20400 -5715
rect 20000 -7295 20020 -5735
rect 20380 -7295 20400 -5735
rect 20000 -7315 20400 -7295
rect 20800 -5735 21200 -5715
rect 20800 -7295 20820 -5735
rect 21180 -7295 21200 -5735
rect 20800 -7315 21200 -7295
rect 21600 -5735 22000 -5715
rect 21600 -7295 21620 -5735
rect 21980 -7295 22000 -5735
rect 21600 -7315 22000 -7295
rect 22400 -5735 22800 -5715
rect 22400 -7295 22420 -5735
rect 22780 -7295 22800 -5735
rect 22400 -7315 22800 -7295
rect 23200 -5735 23600 -5715
rect 23200 -7295 23220 -5735
rect 23580 -7295 23600 -5735
rect 23200 -7315 23600 -7295
<< ndiffc >>
rect -380 25 -20 1585
rect 420 25 780 1585
rect 1220 25 1580 1585
rect 2020 25 2380 1585
rect 2820 25 3180 1585
rect 3620 25 3980 1585
rect 4420 25 4780 1585
rect 5220 25 5580 1585
rect 6020 25 6380 1585
rect 6820 25 7180 1585
rect 7620 25 7980 1585
rect 8420 25 8780 1585
rect 9220 25 9580 1585
rect 10020 25 10380 1585
rect 10820 25 11180 1585
rect 11620 25 11980 1585
rect 12420 25 12780 1585
rect 13220 25 13580 1585
rect 14020 25 14380 1585
rect 14820 25 15180 1585
rect 15620 25 15980 1585
rect 16420 25 16780 1585
rect 18420 25 18780 1585
rect 19220 25 19580 1585
rect 20020 25 20380 1585
rect 20820 25 21180 1585
rect 21620 25 21980 1585
rect 22420 25 22780 1585
rect 23220 25 23580 1585
rect -380 -2375 -20 -815
rect 420 -2375 780 -815
rect 1220 -2375 1580 -815
rect 2020 -2375 2380 -815
rect 2820 -2375 3180 -815
rect 3620 -2375 3980 -815
rect 4420 -2375 4780 -815
rect 5220 -2375 5580 -815
rect 6020 -2375 6380 -815
rect 6820 -2375 7180 -815
rect 7620 -2375 7980 -815
rect 8420 -2375 8780 -815
rect 9220 -2375 9580 -815
rect 10020 -2375 10380 -815
rect 10820 -2375 11180 -815
rect 11620 -2375 11980 -815
rect 12420 -2375 12780 -815
rect 13220 -2375 13580 -815
rect 14020 -2375 14380 -815
rect 14820 -2375 15180 -815
rect 15620 -2375 15980 -815
rect 16420 -2375 16780 -815
rect 18420 -2375 18780 -815
rect 19220 -2375 19580 -815
rect 20020 -2375 20380 -815
rect 20820 -2375 21180 -815
rect 21620 -2375 21980 -815
rect 22420 -2375 22780 -815
rect 23220 -2375 23580 -815
rect -380 -4895 -20 -3335
rect 420 -4895 780 -3335
rect 1220 -4895 1580 -3335
rect 2020 -4895 2380 -3335
rect 2820 -4895 3180 -3335
rect 3620 -4895 3980 -3335
rect 4420 -4895 4780 -3335
rect 5220 -4895 5580 -3335
rect 6020 -4895 6380 -3335
rect 6820 -4895 7180 -3335
rect 7620 -4895 7980 -3335
rect 8420 -4895 8780 -3335
rect 9220 -4895 9580 -3335
rect 10020 -4895 10380 -3335
rect 10820 -4895 11180 -3335
rect 11620 -4895 11980 -3335
rect 12420 -4895 12780 -3335
rect 13220 -4895 13580 -3335
rect 14020 -4895 14380 -3335
rect 14820 -4895 15180 -3335
rect 15620 -4895 15980 -3335
rect 16420 -4895 16780 -3335
rect 18420 -4895 18780 -3335
rect 19220 -4895 19580 -3335
rect 20020 -4895 20380 -3335
rect 20820 -4895 21180 -3335
rect 21620 -4895 21980 -3335
rect 22420 -4895 22780 -3335
rect 23220 -4895 23580 -3335
rect -380 -7295 -20 -5735
rect 420 -7295 780 -5735
rect 1220 -7295 1580 -5735
rect 2020 -7295 2380 -5735
rect 2820 -7295 3180 -5735
rect 3620 -7295 3980 -5735
rect 4420 -7295 4780 -5735
rect 5220 -7295 5580 -5735
rect 6020 -7295 6380 -5735
rect 6820 -7295 7180 -5735
rect 7620 -7295 7980 -5735
rect 8420 -7295 8780 -5735
rect 9220 -7295 9580 -5735
rect 10020 -7295 10380 -5735
rect 10820 -7295 11180 -5735
rect 11620 -7295 11980 -5735
rect 12420 -7295 12780 -5735
rect 13220 -7295 13580 -5735
rect 14015 -7295 14380 -5735
rect 14820 -7295 15180 -5735
rect 15620 -7295 15980 -5735
rect 16420 -7295 16780 -5735
rect 18420 -7295 18780 -5735
rect 19220 -7295 19580 -5735
rect 20020 -7295 20380 -5735
rect 20820 -7295 21180 -5735
rect 21620 -7295 21980 -5735
rect 22420 -7295 22780 -5735
rect 23220 -7295 23580 -5735
<< psubdiff >>
rect 5370 2015 5420 2030
rect 5370 1995 5385 2015
rect 5405 1995 5420 2015
rect 5370 1980 5420 1995
rect 1375 1760 1425 1775
rect 1375 1740 1390 1760
rect 1410 1740 1425 1760
rect 1375 1725 1425 1740
rect 3765 1760 3815 1775
rect 8175 1765 8225 1780
rect 3765 1740 3780 1760
rect 3800 1740 3815 1760
rect 3765 1725 3815 1740
rect 8175 1745 8190 1765
rect 8210 1745 8225 1765
rect 8175 1730 8225 1745
rect 14180 1830 14230 1845
rect 14180 1810 14195 1830
rect 14215 1810 14230 1830
rect 14180 1795 14230 1810
rect -800 1585 -400 1605
rect -800 25 -780 1585
rect -420 25 -400 1585
rect -800 5 -400 25
rect 11200 1585 11600 1605
rect 11200 25 11220 1585
rect 11580 25 11600 1585
rect 11200 5 11600 25
rect 16800 1585 17200 1605
rect 16800 25 16820 1585
rect 17180 25 17200 1585
rect 16800 5 17200 25
rect 18000 1585 18400 1605
rect 18000 25 18020 1585
rect 18380 25 18400 1585
rect 18000 5 18400 25
rect 23600 1585 24000 1605
rect 23600 25 23620 1585
rect 23980 25 24000 1585
rect 23600 5 24000 25
rect 1375 -240 1425 -225
rect 1375 -260 1390 -240
rect 1410 -260 1425 -240
rect 1375 -275 1425 -260
rect 3765 -240 3815 -225
rect 3765 -260 3780 -240
rect 3800 -260 3815 -240
rect 3765 -275 3815 -260
rect 5370 -235 5420 -220
rect 5370 -255 5385 -235
rect 5405 -255 5420 -235
rect 5370 -270 5420 -255
rect 8175 -235 8225 -220
rect 8175 -255 8190 -235
rect 8210 -255 8225 -235
rect 8175 -270 8225 -255
rect 14180 -170 14230 -155
rect 14180 -190 14195 -170
rect 14215 -190 14230 -170
rect 14180 -205 14230 -190
rect -800 -815 -400 -795
rect -800 -2375 -780 -815
rect -420 -2375 -400 -815
rect -800 -2395 -400 -2375
rect 11200 -815 11600 -795
rect 11200 -2375 11220 -815
rect 11580 -2375 11600 -815
rect 11200 -2395 11600 -2375
rect 16800 -815 17200 -795
rect 16800 -2375 16820 -815
rect 17180 -2375 17200 -815
rect 16800 -2395 17200 -2375
rect 18000 -815 18400 -795
rect 18000 -2375 18020 -815
rect 18380 -2375 18400 -815
rect 18000 -2395 18400 -2375
rect 23600 -815 24000 -795
rect 23600 -2375 23620 -815
rect 23980 -2375 24000 -815
rect 23600 -2395 24000 -2375
rect 2175 -2670 2225 -2655
rect 2175 -2690 2190 -2670
rect 2210 -2690 2225 -2670
rect 2175 -2705 2225 -2690
rect 4560 -2670 4610 -2655
rect 4560 -2690 4575 -2670
rect 4595 -2690 4610 -2670
rect 4560 -2705 4610 -2690
rect 6580 -2670 6630 -2655
rect 6580 -2690 6595 -2670
rect 6615 -2690 6630 -2670
rect 6580 -2705 6630 -2690
rect 8580 -2670 8630 -2655
rect 8580 -2690 8595 -2670
rect 8615 -2690 8630 -2670
rect 8580 -2705 8630 -2690
rect 14180 -2670 14230 -2655
rect 14180 -2690 14195 -2670
rect 14215 -2690 14230 -2670
rect 14180 -2705 14230 -2690
rect -800 -3335 -400 -3315
rect -800 -4895 -780 -3335
rect -420 -4895 -400 -3335
rect -800 -4915 -400 -4895
rect 11200 -3335 11600 -3315
rect 11200 -4895 11220 -3335
rect 11580 -4895 11600 -3335
rect 11200 -4915 11600 -4895
rect 16800 -3335 17200 -3315
rect 16800 -4895 16820 -3335
rect 17180 -4895 17200 -3335
rect 16800 -4915 17200 -4895
rect 18000 -3335 18400 -3315
rect 18000 -4895 18020 -3335
rect 18380 -4895 18400 -3335
rect 18000 -4915 18400 -4895
rect 23600 -3335 24000 -3315
rect 23600 -4895 23620 -3335
rect 23980 -4895 24000 -3335
rect 23600 -4915 24000 -4895
rect 2175 -5170 2225 -5155
rect 2175 -5190 2190 -5170
rect 2210 -5190 2225 -5170
rect 2175 -5205 2225 -5190
rect 4560 -5170 4610 -5155
rect 4560 -5190 4575 -5170
rect 4595 -5190 4610 -5170
rect 4560 -5205 4610 -5190
rect 6580 -5170 6630 -5155
rect 6580 -5190 6595 -5170
rect 6615 -5190 6630 -5170
rect 6580 -5205 6630 -5190
rect 8580 -5170 8630 -5155
rect 8580 -5190 8595 -5170
rect 8615 -5190 8630 -5170
rect 8580 -5205 8630 -5190
rect 10580 -5170 10630 -5155
rect 10580 -5190 10595 -5170
rect 10615 -5190 10630 -5170
rect 10580 -5205 10630 -5190
rect 14180 -5170 14230 -5155
rect 14180 -5190 14195 -5170
rect 14215 -5190 14230 -5170
rect 14180 -5205 14230 -5190
rect -800 -5735 -400 -5715
rect -800 -7295 -780 -5735
rect -420 -7295 -400 -5735
rect -800 -7315 -400 -7295
rect 11200 -5735 11600 -5715
rect 11200 -7295 11220 -5735
rect 11580 -7295 11600 -5735
rect 11200 -7315 11600 -7295
rect 16800 -5735 17200 -5715
rect 16800 -7295 16820 -5735
rect 17180 -7295 17200 -5735
rect 16800 -7315 17200 -7295
rect 18000 -5735 18400 -5715
rect 18000 -7295 18020 -5735
rect 18380 -7295 18400 -5735
rect 18000 -7315 18400 -7295
rect 23600 -5735 24000 -5715
rect 23600 -7295 23620 -5735
rect 23980 -7295 24000 -5735
rect 23600 -7315 24000 -7295
rect 2175 -7370 2225 -7355
rect 2175 -7390 2190 -7370
rect 2210 -7390 2225 -7370
rect 2175 -7405 2225 -7390
rect 4575 -7360 4625 -7345
rect 4575 -7380 4590 -7360
rect 4610 -7380 4625 -7360
rect 4575 -7395 4625 -7380
rect 6175 -7370 6225 -7355
rect 6175 -7390 6190 -7370
rect 6210 -7390 6225 -7370
rect 6175 -7405 6225 -7390
rect 8575 -7360 8625 -7345
rect 8575 -7380 8590 -7360
rect 8610 -7380 8625 -7360
rect 8575 -7395 8625 -7380
rect 14180 -7360 14230 -7345
rect 14180 -7380 14195 -7360
rect 14215 -7380 14230 -7360
rect 14180 -7395 14230 -7380
<< psubdiffcont >>
rect 5385 1995 5405 2015
rect 1390 1740 1410 1760
rect 3780 1740 3800 1760
rect 8190 1745 8210 1765
rect 14195 1810 14215 1830
rect -780 25 -420 1585
rect 11220 25 11580 1585
rect 16820 25 17180 1585
rect 18020 25 18380 1585
rect 23620 25 23980 1585
rect 1390 -260 1410 -240
rect 3780 -260 3800 -240
rect 5385 -255 5405 -235
rect 8190 -255 8210 -235
rect 14195 -190 14215 -170
rect -780 -2375 -420 -815
rect 11220 -2375 11580 -815
rect 16820 -2375 17180 -815
rect 18020 -2375 18380 -815
rect 23620 -2375 23980 -815
rect 2190 -2690 2210 -2670
rect 4575 -2690 4595 -2670
rect 6595 -2690 6615 -2670
rect 8595 -2690 8615 -2670
rect 14195 -2690 14215 -2670
rect -780 -4895 -420 -3335
rect 11220 -4895 11580 -3335
rect 16820 -4895 17180 -3335
rect 18020 -4895 18380 -3335
rect 23620 -4895 23980 -3335
rect 2190 -5190 2210 -5170
rect 4575 -5190 4595 -5170
rect 6595 -5190 6615 -5170
rect 8595 -5190 8615 -5170
rect 10595 -5190 10615 -5170
rect 14195 -5190 14215 -5170
rect -780 -7295 -420 -5735
rect 11220 -7295 11580 -5735
rect 16820 -7295 17180 -5735
rect 18020 -7295 18380 -5735
rect 23620 -7295 23980 -5735
rect 2190 -7390 2210 -7370
rect 4590 -7380 4610 -7360
rect 6190 -7390 6210 -7370
rect 8590 -7380 8610 -7360
rect 14195 -7380 14215 -7360
<< poly >>
rect 4000 1725 6800 1765
rect 3200 1710 3600 1720
rect 3200 1630 3220 1710
rect 3580 1630 3600 1710
rect 0 1605 400 1620
rect 800 1605 1200 1620
rect 1600 1605 2000 1620
rect 2400 1605 2800 1620
rect 3200 1605 3600 1630
rect 4000 1605 4400 1725
rect 4800 1605 5200 1725
rect 5600 1605 6000 1725
rect 6400 1605 6800 1725
rect 7200 1710 7600 1720
rect 7200 1630 7220 1710
rect 7580 1630 7600 1710
rect 7200 1605 7600 1630
rect 8000 1605 8400 1620
rect 8800 1605 9200 1925
rect 9600 1605 10000 1620
rect 10400 1605 10800 1620
rect 12000 1605 12400 1620
rect 12800 1605 13200 1620
rect 13600 1605 14000 1620
rect 14400 1605 14800 1620
rect 15200 1605 15600 1620
rect 16000 1605 16400 1620
rect 18800 1605 19200 1620
rect 19600 1605 20000 1620
rect 20400 1605 20800 1620
rect 21200 1605 21600 1620
rect 22000 1605 22400 1620
rect 22800 1605 23200 1620
rect 0 -10 400 5
rect 800 -10 1200 5
rect -390 -20 1200 -10
rect -390 -100 -380 -20
rect -20 -100 420 -20
rect 780 -100 1200 -20
rect -390 -110 1200 -100
rect 1600 -115 2000 5
rect 2400 -115 2800 5
rect 3200 -10 3600 5
rect 4000 -10 4400 5
rect 4800 -10 5200 5
rect 5600 -10 6000 5
rect 6400 -10 6800 5
rect 7200 -10 7600 5
rect 5950 -20 5990 -10
rect 5950 -40 5960 -20
rect 5980 -40 5990 -20
rect 5950 -50 5990 -40
rect 6410 -20 6450 -10
rect 6410 -40 6420 -20
rect 6440 -40 6450 -20
rect 6410 -50 6450 -40
rect 8000 -115 8400 5
rect 8800 -115 9200 5
rect 9600 -10 10000 5
rect 10400 -10 10800 5
rect 12000 -10 12400 5
rect 9600 -20 11190 -10
rect 9600 -100 10020 -20
rect 10380 -100 10820 -20
rect 11180 -100 11190 -20
rect 9600 -110 11190 -100
rect 11610 -20 12400 -10
rect 11610 -100 11620 -20
rect 11980 -100 12400 -20
rect 11610 -110 12400 -100
rect 1600 -120 9200 -115
rect 1600 -150 6815 -120
rect 7185 -150 9200 -120
rect 1600 -155 9200 -150
rect 3200 -690 3600 -680
rect 3200 -770 3220 -690
rect 3580 -770 3600 -690
rect 7200 -690 7600 -680
rect 0 -795 400 -780
rect 800 -795 1200 -780
rect 1600 -795 2000 -780
rect 2400 -795 2800 -780
rect 3200 -795 3600 -770
rect 5950 -750 5990 -740
rect 5950 -770 5960 -750
rect 5980 -770 5990 -750
rect 5950 -780 5990 -770
rect 6410 -750 6450 -740
rect 6410 -770 6420 -750
rect 6440 -770 6450 -750
rect 6410 -780 6450 -770
rect 7200 -770 7220 -690
rect 7580 -770 7600 -690
rect 12800 -715 13200 5
rect 13600 -715 14000 5
rect 14400 -715 14800 5
rect 15200 -715 15600 5
rect 16000 -10 16400 5
rect 18800 -10 19200 5
rect 16000 -20 16790 -10
rect 16000 -100 16420 -20
rect 16780 -100 16790 -20
rect 16000 -110 16790 -100
rect 18410 -20 19200 -10
rect 18410 -100 18420 -20
rect 18780 -100 19200 -20
rect 18410 -110 19200 -100
rect 12750 -725 15600 -715
rect 12750 -745 12760 -725
rect 12780 -745 15600 -725
rect 12750 -755 15600 -745
rect 4000 -795 4400 -780
rect 4800 -795 5200 -780
rect 5600 -795 6000 -780
rect 6400 -795 6800 -780
rect 7200 -795 7600 -770
rect 8000 -795 8400 -780
rect 8800 -795 9200 -780
rect 9600 -795 10000 -780
rect 10400 -795 10800 -780
rect 12000 -795 12400 -780
rect 12800 -795 13200 -755
rect 13600 -795 14000 -755
rect 14400 -795 14800 -755
rect 15200 -795 15600 -755
rect 16000 -795 16400 -780
rect 18800 -795 19200 -780
rect 19600 -795 20000 5
rect 20400 -795 20800 5
rect 21200 -795 21600 5
rect 22000 -795 22400 5
rect 22800 -10 23200 5
rect 22800 -20 23590 -10
rect 22800 -100 23220 -20
rect 23580 -100 23590 -20
rect 22800 -110 23590 -100
rect 22800 -795 23200 -780
rect 0 -2410 400 -2395
rect 800 -2410 1200 -2395
rect -390 -2420 1200 -2410
rect -390 -2500 -380 -2420
rect -20 -2500 420 -2420
rect 780 -2500 1200 -2420
rect -390 -2510 1200 -2500
rect 1600 -2515 2000 -2395
rect 2400 -2515 2800 -2395
rect 3200 -2410 3600 -2395
rect 4000 -2450 4400 -2395
rect 4800 -2450 5200 -2395
rect 5600 -2450 6000 -2395
rect 6400 -2450 6800 -2395
rect 7200 -2410 7600 -2395
rect 4000 -2490 6800 -2450
rect 8000 -2515 8400 -2395
rect 8800 -2515 9200 -2395
rect 9600 -2410 10000 -2395
rect 10400 -2410 10800 -2395
rect 12000 -2410 12400 -2395
rect 12800 -2410 13200 -2395
rect 13600 -2410 14000 -2395
rect 14400 -2410 14800 -2395
rect 15200 -2410 15600 -2395
rect 16000 -2410 16400 -2395
rect 18800 -2410 19200 -2395
rect 9600 -2420 11190 -2410
rect 9600 -2500 10020 -2420
rect 10380 -2500 10820 -2420
rect 11180 -2500 11190 -2420
rect 9600 -2510 11190 -2500
rect 11610 -2420 12400 -2410
rect 11610 -2500 11620 -2420
rect 11980 -2500 12400 -2420
rect 11610 -2510 12400 -2500
rect 16000 -2420 16790 -2410
rect 16000 -2500 16420 -2420
rect 16780 -2500 16790 -2420
rect 16000 -2510 16790 -2500
rect 18410 -2420 19200 -2410
rect 18410 -2500 18420 -2420
rect 18780 -2500 19200 -2420
rect 18410 -2510 19200 -2500
rect 1600 -2555 9200 -2515
rect 7200 -3270 7600 -3260
rect 7200 -3290 7570 -3270
rect 7590 -3290 7600 -3270
rect 0 -3315 400 -3300
rect 800 -3315 1200 -3300
rect 1600 -3315 2000 -3300
rect 2400 -3315 2800 -3300
rect 3200 -3315 3600 -3300
rect 4000 -3315 4400 -3300
rect 4800 -3315 5200 -3300
rect 5600 -3315 6000 -3300
rect 6400 -3315 6800 -3300
rect 7200 -3315 7600 -3290
rect 8000 -3315 8400 -3300
rect 8800 -3315 9200 -3300
rect 9600 -3315 10000 -3300
rect 10400 -3315 10800 -3300
rect 12000 -3315 12400 -3300
rect 12800 -3315 13200 -3300
rect 13600 -3315 14000 -3300
rect 14400 -3315 14800 -3300
rect 15200 -3315 15600 -3300
rect 16000 -3315 16400 -3300
rect 18800 -3315 19200 -3300
rect 19600 -3315 20000 -2395
rect 20400 -3315 20800 -2395
rect 21200 -3315 21600 -2395
rect 22000 -3315 22400 -2395
rect 22800 -2410 23200 -2395
rect 22800 -2420 23590 -2410
rect 22800 -2500 23220 -2420
rect 23580 -2500 23590 -2420
rect 22800 -2510 23590 -2500
rect 22800 -3315 23200 -3300
rect 0 -4930 400 -4915
rect -390 -4940 400 -4930
rect -390 -5020 -380 -4940
rect -20 -5020 400 -4940
rect -390 -5030 400 -5020
rect 800 -4955 1200 -4915
rect 800 -4965 1250 -4955
rect 800 -4985 1220 -4965
rect 1240 -4985 1250 -4965
rect 800 -4995 1250 -4985
rect 1600 -4995 2000 -4915
rect 2400 -4955 2800 -4915
rect 2400 -4965 2850 -4955
rect 2400 -4985 2820 -4965
rect 2840 -4985 2850 -4965
rect 2400 -4995 2850 -4985
rect 3200 -4995 3600 -4915
rect 4000 -4930 4400 -4915
rect 4000 -4940 4450 -4930
rect 4000 -4960 4420 -4940
rect 4440 -4960 4450 -4940
rect 4000 -4970 4450 -4960
rect 4800 -4995 5200 -4915
rect 5600 -4995 6000 -4915
rect 6400 -4930 6800 -4915
rect 6585 -4940 6625 -4930
rect 6585 -4960 6595 -4940
rect 6615 -4960 6625 -4940
rect 6585 -4970 6625 -4960
rect 800 -5025 6000 -4995
rect 800 -5605 1200 -5025
rect 1600 -5605 2000 -5025
rect 2400 -5605 2800 -5025
rect 3200 -5605 3600 -5025
rect 4800 -5605 5200 -5025
rect 5600 -5605 6000 -5025
rect 7200 -4995 7600 -4915
rect 8000 -4995 8400 -4915
rect 8800 -4995 9200 -4915
rect 9600 -4995 10000 -4915
rect 7200 -5025 10000 -4995
rect 800 -5635 6000 -5605
rect 800 -5645 1250 -5635
rect 800 -5665 1220 -5645
rect 1240 -5665 1250 -5645
rect 800 -5675 1250 -5665
rect 1600 -5645 2050 -5635
rect 1600 -5665 2020 -5645
rect 2040 -5665 2050 -5645
rect 1600 -5675 2050 -5665
rect 2400 -5645 2850 -5635
rect 2400 -5665 2820 -5645
rect 2840 -5665 2850 -5645
rect 2400 -5675 2850 -5665
rect 0 -5715 400 -5700
rect 800 -5715 1200 -5675
rect 1600 -5715 2000 -5675
rect 2400 -5715 2800 -5675
rect 3200 -5715 3600 -5635
rect 4000 -5670 4450 -5660
rect 4000 -5690 4420 -5670
rect 4440 -5690 4450 -5670
rect 4000 -5700 4450 -5690
rect 4000 -5715 4400 -5700
rect 4800 -5715 5200 -5635
rect 5600 -5715 6000 -5635
rect 7200 -5605 7600 -5025
rect 8000 -5605 8400 -5025
rect 8800 -5605 9200 -5025
rect 9600 -5605 10000 -5025
rect 10400 -4930 10800 -4915
rect 12000 -4930 12400 -4915
rect 10400 -4940 11190 -4930
rect 10400 -5020 10820 -4940
rect 11180 -5020 11190 -4940
rect 10400 -5030 11190 -5020
rect 11610 -4940 12400 -4930
rect 11610 -5020 11620 -4940
rect 11980 -5020 12400 -4940
rect 11610 -5030 12400 -5020
rect 12800 -5605 13200 -4915
rect 7200 -5635 13200 -5605
rect 6585 -5670 6625 -5660
rect 6585 -5690 6595 -5670
rect 6615 -5690 6625 -5670
rect 6585 -5700 6625 -5690
rect 6400 -5715 6800 -5700
rect 7200 -5715 7600 -5635
rect 8000 -5715 8400 -5635
rect 8800 -5715 9200 -5635
rect 9600 -5645 10050 -5635
rect 9600 -5665 10020 -5645
rect 10040 -5665 10050 -5645
rect 9600 -5675 10050 -5665
rect 9600 -5715 10000 -5675
rect 10400 -5715 10800 -5700
rect 12000 -5715 12400 -5700
rect 12800 -5715 13200 -5635
rect 13600 -5715 14000 -4915
rect 14400 -5605 14800 -4915
rect 15200 -5605 15600 -4915
rect 16000 -4930 16400 -4915
rect 18800 -4930 19200 -4915
rect 19600 -4930 20000 -4915
rect 20400 -4930 20800 -4915
rect 21200 -4930 21600 -4915
rect 22000 -4930 22400 -4915
rect 22800 -4930 23200 -4915
rect 16000 -4940 16790 -4930
rect 16000 -5020 16420 -4940
rect 16780 -5020 16790 -4940
rect 16000 -5030 16790 -5020
rect 18410 -4940 19200 -4930
rect 18410 -5020 18420 -4940
rect 18780 -5020 19200 -4940
rect 18410 -5030 19200 -5020
rect 22800 -4940 23590 -4930
rect 22800 -5020 23220 -4940
rect 23580 -5020 23590 -4940
rect 22800 -5030 23590 -5020
rect 14400 -5645 17635 -5605
rect 14400 -5715 14800 -5645
rect 15200 -5715 15600 -5645
rect 16000 -5715 16400 -5700
rect 18800 -5715 19200 -5700
rect 19600 -5715 20000 -5700
rect 20400 -5715 20800 -5700
rect 21200 -5715 21600 -5700
rect 22000 -5715 22400 -5700
rect 22800 -5715 23200 -5700
rect 0 -7330 400 -7315
rect 800 -7330 1200 -7315
rect 1600 -7330 2000 -7315
rect 2400 -7330 2800 -7315
rect 3200 -7330 3600 -7315
rect 4000 -7330 4400 -7315
rect 4800 -7330 5200 -7315
rect 5600 -7330 6000 -7315
rect 6400 -7330 6800 -7315
rect -390 -7340 400 -7330
rect -390 -7420 -380 -7340
rect -20 -7420 400 -7340
rect 7200 -7340 7600 -7315
rect -390 -7430 400 -7420
rect 7200 -7420 7210 -7340
rect 7590 -7420 7600 -7340
rect 7200 -7430 7600 -7420
rect 8000 -7340 8400 -7315
rect 8000 -7420 8010 -7340
rect 8390 -7420 8400 -7340
rect 8800 -7340 9200 -7315
rect 8000 -7430 8400 -7420
rect 8800 -7420 8810 -7340
rect 9190 -7420 9200 -7340
rect 8800 -7430 9200 -7420
rect 9600 -7340 10000 -7315
rect 9600 -7420 9610 -7340
rect 9990 -7420 10000 -7340
rect 9600 -7430 10000 -7420
rect 10400 -7330 10800 -7315
rect 12000 -7330 12400 -7315
rect 10400 -7340 11190 -7330
rect 10400 -7420 10820 -7340
rect 11180 -7420 11190 -7340
rect 10400 -7430 11190 -7420
rect 11610 -7340 12400 -7330
rect 11610 -7420 11620 -7340
rect 11980 -7420 12400 -7340
rect 11610 -7430 12400 -7420
rect 12800 -7340 13200 -7315
rect 12800 -7420 12810 -7340
rect 13190 -7420 13200 -7340
rect 12800 -7430 13200 -7420
rect 13600 -7340 14000 -7315
rect 14400 -7330 14800 -7315
rect 15200 -7330 15600 -7315
rect 16000 -7330 16400 -7315
rect 18800 -7330 19200 -7315
rect 13600 -7420 13610 -7340
rect 13990 -7420 14000 -7340
rect 16000 -7340 16790 -7330
rect 13600 -7430 14000 -7420
rect 16000 -7420 16420 -7340
rect 16780 -7420 16790 -7340
rect 16000 -7430 16790 -7420
rect 18410 -7340 19200 -7330
rect 18410 -7420 18420 -7340
rect 18780 -7420 19200 -7340
rect 18410 -7430 19200 -7420
rect 19600 -7340 20000 -7315
rect 19600 -7420 19610 -7340
rect 19990 -7420 20000 -7340
rect 19600 -7430 20000 -7420
rect 20400 -7340 20800 -7315
rect 20400 -7420 20410 -7340
rect 20790 -7420 20800 -7340
rect 20400 -7430 20800 -7420
rect 21200 -7340 21600 -7315
rect 21200 -7420 21210 -7340
rect 21590 -7420 21600 -7340
rect 21200 -7430 21600 -7420
rect 22000 -7340 22400 -7315
rect 22000 -7420 22010 -7340
rect 22390 -7420 22400 -7340
rect 22000 -7430 22400 -7420
rect 22800 -7330 23200 -7315
rect 22800 -7340 23590 -7330
rect 22800 -7420 23220 -7340
rect 23580 -7420 23590 -7340
rect 22800 -7430 23590 -7420
<< polycont >>
rect 3220 1630 3580 1710
rect 7220 1630 7580 1710
rect -380 -100 -20 -20
rect 420 -100 780 -20
rect 5960 -40 5980 -20
rect 6420 -40 6440 -20
rect 10020 -100 10380 -20
rect 10820 -100 11180 -20
rect 11620 -100 11980 -20
rect 6815 -150 7185 -120
rect 3220 -770 3580 -690
rect 5960 -770 5980 -750
rect 6420 -770 6440 -750
rect 7220 -770 7580 -690
rect 16420 -100 16780 -20
rect 18420 -100 18780 -20
rect 12760 -745 12780 -725
rect 23220 -100 23580 -20
rect -380 -2500 -20 -2420
rect 420 -2500 780 -2420
rect 10020 -2500 10380 -2420
rect 10820 -2500 11180 -2420
rect 11620 -2500 11980 -2420
rect 16420 -2500 16780 -2420
rect 18420 -2500 18780 -2420
rect 7570 -3290 7590 -3270
rect 23220 -2500 23580 -2420
rect -380 -5020 -20 -4940
rect 1220 -4985 1240 -4965
rect 2820 -4985 2840 -4965
rect 4420 -4960 4440 -4940
rect 6595 -4960 6615 -4940
rect 1220 -5665 1240 -5645
rect 2020 -5665 2040 -5645
rect 2820 -5665 2840 -5645
rect 4420 -5690 4440 -5670
rect 10820 -5020 11180 -4940
rect 11620 -5020 11980 -4940
rect 6595 -5690 6615 -5670
rect 10020 -5665 10040 -5645
rect 16420 -5020 16780 -4940
rect 18420 -5020 18780 -4940
rect 23220 -5020 23580 -4940
rect -380 -7420 -20 -7340
rect 7210 -7420 7590 -7340
rect 8010 -7420 8390 -7340
rect 8810 -7420 9190 -7340
rect 9610 -7420 9990 -7340
rect 10820 -7420 11180 -7340
rect 11620 -7420 11980 -7340
rect 12810 -7420 13190 -7340
rect 13610 -7420 13990 -7340
rect 16420 -7420 16780 -7340
rect 18420 -7420 18780 -7340
rect 19610 -7420 19990 -7340
rect 20410 -7420 20790 -7340
rect 21210 -7420 21590 -7340
rect 22010 -7420 22390 -7340
rect 23220 -7420 23580 -7340
<< locali >>
rect 5375 2060 5415 2070
rect 5375 2040 5385 2060
rect 5405 2040 5415 2060
rect 5375 2015 5415 2040
rect 5375 1995 5385 2015
rect 5405 1995 5415 2015
rect 5375 1985 5415 1995
rect 14185 1875 14225 1885
rect 14185 1855 14195 1875
rect 14215 1855 14225 1875
rect 14185 1830 14225 1855
rect 3200 1820 3600 1830
rect 1380 1805 1420 1815
rect 1380 1785 1390 1805
rect 1410 1785 1420 1805
rect 1380 1760 1420 1785
rect 1380 1740 1390 1760
rect 1410 1740 1420 1760
rect 1380 1730 1420 1740
rect 3200 1730 3210 1820
rect 3590 1730 3600 1820
rect 3770 1805 3810 1815
rect 3770 1785 3780 1805
rect 3800 1785 3810 1805
rect 3770 1760 3810 1785
rect 3770 1740 3780 1760
rect 3800 1740 3810 1760
rect 3770 1730 3810 1740
rect 8180 1810 8220 1820
rect 8180 1790 8190 1810
rect 8210 1790 8220 1810
rect 14185 1810 14195 1830
rect 14215 1810 14225 1830
rect 14185 1800 14225 1810
rect 8180 1765 8220 1790
rect 8180 1745 8190 1765
rect 8210 1745 8220 1765
rect 8180 1735 8220 1745
rect 3200 1720 3600 1730
rect 3210 1710 3590 1720
rect 3210 1630 3220 1710
rect 3580 1630 3590 1710
rect 3210 1620 3590 1630
rect 7210 1710 7590 1720
rect 7210 1630 7220 1710
rect 7580 1630 7590 1710
rect 7210 1620 7590 1630
rect 20200 1645 21800 1745
rect 20200 1595 20390 1645
rect 21610 1595 21800 1645
rect -790 1585 -10 1595
rect -790 25 -780 1585
rect -420 25 -380 1585
rect -20 25 -10 1585
rect -790 15 -10 25
rect -390 -20 -10 15
rect -390 -100 -380 -20
rect -20 -100 -10 -20
rect -390 -110 -10 -100
rect 410 1585 790 1595
rect 410 25 420 1585
rect 780 25 790 1585
rect 410 -20 790 25
rect 1210 1585 1590 1595
rect 1210 25 1220 1585
rect 1580 25 1590 1585
rect 1210 15 1590 25
rect 2010 1585 2390 1595
rect 2010 25 2020 1585
rect 2380 25 2390 1585
rect 410 -100 420 -20
rect 780 -100 790 -20
rect 410 -110 790 -100
rect 1380 -195 1420 -185
rect 1380 -215 1390 -195
rect 1410 -215 1420 -195
rect 1380 -240 1420 -215
rect 1380 -260 1390 -240
rect 1410 -260 1420 -240
rect 1380 -270 1420 -260
rect -790 -815 -10 -805
rect -790 -2375 -780 -815
rect -420 -2375 -380 -815
rect -20 -2375 -10 -815
rect -790 -2385 -10 -2375
rect -390 -2420 -10 -2385
rect -390 -2500 -380 -2420
rect -20 -2500 -10 -2420
rect -390 -2510 -10 -2500
rect 410 -815 790 -805
rect 410 -2375 420 -815
rect 780 -2375 790 -815
rect 410 -2420 790 -2375
rect 1210 -815 1590 -805
rect 1210 -2375 1220 -815
rect 1580 -2375 1590 -815
rect 1210 -2385 1590 -2375
rect 2010 -815 2390 25
rect 2810 1585 3190 1595
rect 2810 25 2820 1585
rect 3180 25 3190 1585
rect 2810 15 3190 25
rect 3610 1585 3990 1595
rect 3610 25 3620 1585
rect 3980 25 3990 1585
rect 3610 15 3990 25
rect 4410 1585 4790 1595
rect 4410 25 4420 1585
rect 4780 25 4790 1585
rect 3770 -195 3810 -185
rect 3770 -215 3780 -195
rect 3800 -215 3810 -195
rect 3770 -240 3810 -215
rect 3770 -260 3780 -240
rect 3800 -260 3810 -240
rect 3770 -270 3810 -260
rect 3200 -575 3600 -565
rect 3200 -670 3210 -575
rect 3590 -670 3600 -575
rect 3200 -680 3600 -670
rect 3210 -690 3590 -680
rect 3210 -770 3220 -690
rect 3580 -770 3590 -690
rect 3210 -780 3590 -770
rect 2010 -2375 2020 -815
rect 2380 -2375 2390 -815
rect 2010 -2385 2390 -2375
rect 2810 -815 3190 -805
rect 2810 -2375 2820 -815
rect 3180 -2375 3190 -815
rect 410 -2500 420 -2420
rect 780 -2500 790 -2420
rect 410 -2510 790 -2500
rect 2180 -2625 2220 -2615
rect 2180 -2645 2190 -2625
rect 2210 -2645 2220 -2625
rect 2180 -2670 2220 -2645
rect 2180 -2690 2190 -2670
rect 2210 -2690 2220 -2670
rect 2180 -2700 2220 -2690
rect -790 -3335 -10 -3325
rect -790 -4895 -780 -3335
rect -420 -4895 -380 -3335
rect -20 -4895 -10 -3335
rect -790 -4905 -10 -4895
rect -390 -4940 -10 -4905
rect -390 -5020 -380 -4940
rect -20 -5020 -10 -4940
rect -390 -5030 -10 -5020
rect 410 -3335 790 -3325
rect 410 -4895 420 -3335
rect 780 -4895 790 -3335
rect 410 -5055 790 -4895
rect 1210 -3335 1590 -3325
rect 1210 -4895 1220 -3335
rect 1580 -4895 1590 -3335
rect 1210 -4955 1590 -4895
rect 2010 -3335 2390 -3325
rect 2010 -4895 2020 -3335
rect 2380 -4895 2390 -3335
rect 1210 -4965 1250 -4955
rect 1210 -4985 1220 -4965
rect 1240 -4985 1250 -4965
rect 1210 -4995 1250 -4985
rect 2010 -5055 2390 -4895
rect 2810 -3335 3190 -2375
rect 3610 -815 3990 -805
rect 3610 -2375 3620 -815
rect 3980 -2375 3990 -815
rect 3610 -2385 3990 -2375
rect 4410 -815 4790 25
rect 5210 1585 5590 1595
rect 5210 25 5220 1585
rect 5580 25 5590 1585
rect 5210 15 5590 25
rect 6010 1585 6390 1595
rect 6010 25 6020 1585
rect 6380 25 6390 1585
rect 5950 -20 5990 -10
rect 5950 -40 5960 -20
rect 5980 -40 5990 -20
rect 5950 -60 5990 -40
rect 5950 -80 5960 -60
rect 5980 -80 5990 -60
rect 5950 -90 5990 -80
rect 5375 -190 5415 -180
rect 5375 -210 5385 -190
rect 5405 -210 5415 -190
rect 5375 -235 5415 -210
rect 5375 -255 5385 -235
rect 5405 -255 5415 -235
rect 5375 -265 5415 -255
rect 5950 -710 5990 -700
rect 5950 -730 5960 -710
rect 5980 -730 5990 -710
rect 5950 -750 5990 -730
rect 5950 -770 5960 -750
rect 5980 -770 5990 -750
rect 5950 -780 5990 -770
rect 4410 -2375 4420 -815
rect 4780 -2375 4790 -815
rect 4410 -2385 4790 -2375
rect 5210 -815 5590 -805
rect 5210 -2375 5220 -815
rect 5580 -2375 5590 -815
rect 5210 -2385 5590 -2375
rect 6010 -815 6390 25
rect 6810 1585 7190 1595
rect 6810 25 6820 1585
rect 7180 25 7190 1585
rect 6410 -20 6450 -10
rect 6410 -40 6420 -20
rect 6440 -40 6450 -20
rect 6410 -60 6450 -40
rect 6410 -80 6420 -60
rect 6440 -80 6450 -60
rect 6410 -90 6450 -80
rect 6810 -120 7190 25
rect 6810 -150 6815 -120
rect 7185 -150 7190 -120
rect 6410 -710 6450 -700
rect 6410 -730 6420 -710
rect 6440 -730 6450 -710
rect 6410 -750 6450 -730
rect 6410 -770 6420 -750
rect 6440 -770 6450 -750
rect 6410 -780 6450 -770
rect 6010 -2375 6020 -815
rect 6380 -2375 6390 -815
rect 6010 -2385 6390 -2375
rect 6810 -815 7190 -150
rect 7610 1585 7990 1595
rect 7610 25 7620 1585
rect 7980 25 7990 1585
rect 7210 -575 7590 -565
rect 7210 -670 7220 -575
rect 7580 -670 7590 -575
rect 7210 -690 7590 -670
rect 7210 -770 7220 -690
rect 7580 -770 7590 -690
rect 7210 -780 7590 -770
rect 6810 -2375 6820 -815
rect 7180 -2375 7190 -815
rect 4565 -2625 4605 -2615
rect 4565 -2645 4575 -2625
rect 4595 -2645 4605 -2625
rect 4565 -2670 4605 -2645
rect 4565 -2690 4575 -2670
rect 4595 -2690 4605 -2670
rect 4565 -2700 4605 -2690
rect 6585 -2625 6625 -2615
rect 6585 -2645 6595 -2625
rect 6615 -2645 6625 -2625
rect 6585 -2670 6625 -2645
rect 6585 -2690 6595 -2670
rect 6615 -2690 6625 -2670
rect 6585 -2700 6625 -2690
rect 6010 -3185 6390 -3175
rect 6010 -3265 6020 -3185
rect 6380 -3265 6390 -3185
rect 2810 -4895 2820 -3335
rect 3180 -4895 3190 -3335
rect 2810 -4955 3190 -4895
rect 3610 -3335 3990 -3325
rect 3610 -4895 3620 -3335
rect 3980 -4895 3990 -3335
rect 2810 -4965 2850 -4955
rect 2810 -4985 2820 -4965
rect 2840 -4985 2850 -4965
rect 2810 -4995 2850 -4985
rect 3610 -5055 3990 -4895
rect 4410 -3335 4790 -3325
rect 4410 -4895 4420 -3335
rect 4780 -4895 4790 -3335
rect 4410 -4930 4790 -4895
rect 5210 -3335 5590 -3325
rect 5210 -4895 5220 -3335
rect 5580 -4895 5590 -3335
rect 4410 -4940 4450 -4930
rect 4410 -4960 4420 -4940
rect 4440 -4960 4450 -4940
rect 4410 -4970 4450 -4960
rect -800 -5095 3990 -5055
rect -790 -5735 -10 -5725
rect -790 -7295 -780 -5735
rect -420 -7295 -380 -5735
rect -20 -7295 -10 -5735
rect -790 -7305 -10 -7295
rect 410 -5735 790 -5095
rect 2180 -5125 2220 -5115
rect 2180 -5145 2190 -5125
rect 2210 -5145 2220 -5125
rect 2180 -5170 2220 -5145
rect 2180 -5190 2190 -5170
rect 2210 -5190 2220 -5170
rect 2180 -5200 2220 -5190
rect 410 -7295 420 -5735
rect 780 -7295 790 -5735
rect 410 -7305 790 -7295
rect 1210 -5645 1250 -5635
rect 1210 -5665 1220 -5645
rect 1240 -5665 1250 -5645
rect 1210 -5675 1250 -5665
rect 2010 -5645 2050 -5635
rect 2010 -5665 2020 -5645
rect 2040 -5665 2050 -5645
rect 2010 -5675 2050 -5665
rect 2810 -5645 2850 -5635
rect 2810 -5665 2820 -5645
rect 2840 -5665 2850 -5645
rect 2810 -5675 2850 -5665
rect 1210 -5735 1590 -5675
rect 1210 -7295 1220 -5735
rect 1580 -7295 1590 -5735
rect 1210 -7305 1590 -7295
rect 2010 -5735 2390 -5675
rect 2010 -7295 2020 -5735
rect 2380 -7295 2390 -5735
rect 2010 -7305 2390 -7295
rect 2810 -5735 3190 -5675
rect 2810 -7295 2820 -5735
rect 3180 -7295 3190 -5735
rect 2810 -7305 3190 -7295
rect 3610 -5735 3990 -5095
rect 4565 -5125 4605 -5115
rect 4565 -5145 4575 -5125
rect 4595 -5145 4605 -5125
rect 4565 -5170 4605 -5145
rect 4565 -5190 4575 -5170
rect 4595 -5190 4605 -5170
rect 4565 -5200 4605 -5190
rect 3610 -7295 3620 -5735
rect 3980 -7295 3990 -5735
rect 3610 -7305 3990 -7295
rect 4410 -5670 4450 -5660
rect 4410 -5690 4420 -5670
rect 4440 -5690 4450 -5670
rect 4410 -5700 4450 -5690
rect 4410 -5735 4790 -5700
rect 4410 -7295 4420 -5735
rect 4780 -7295 4790 -5735
rect 4410 -7305 4790 -7295
rect 5210 -5735 5590 -4895
rect 5210 -7295 5220 -5735
rect 5580 -7295 5590 -5735
rect 5210 -7305 5590 -7295
rect 6010 -3335 6390 -3265
rect 6010 -4895 6020 -3335
rect 6380 -4895 6390 -3335
rect 6010 -5735 6390 -4895
rect 6810 -3335 7190 -2375
rect 7610 -815 7990 25
rect 8410 1585 8790 1595
rect 8410 25 8420 1585
rect 8780 25 8790 1585
rect 8180 -190 8220 -180
rect 8180 -210 8190 -190
rect 8210 -210 8220 -190
rect 8180 -235 8220 -210
rect 8180 -255 8190 -235
rect 8210 -255 8220 -235
rect 8180 -265 8220 -255
rect 7610 -2375 7620 -815
rect 7980 -2375 7990 -815
rect 7610 -3260 7990 -2375
rect 8410 -815 8790 25
rect 9210 1585 9590 1595
rect 9210 25 9220 1585
rect 9580 25 9590 1585
rect 9210 15 9590 25
rect 10010 1585 10390 1595
rect 10010 25 10020 1585
rect 10380 25 10390 1585
rect 10010 -20 10390 25
rect 10010 -100 10020 -20
rect 10380 -100 10390 -20
rect 10010 -110 10390 -100
rect 10810 1585 11990 1595
rect 10810 25 10820 1585
rect 11180 25 11220 1585
rect 11580 25 11620 1585
rect 11980 25 11990 1585
rect 10810 15 11990 25
rect 10810 -20 11190 15
rect 10810 -100 10820 -20
rect 11180 -100 11190 -20
rect 10810 -110 11190 -100
rect 11610 -20 11990 15
rect 11610 -100 11620 -20
rect 11980 -100 11990 -20
rect 11610 -110 11990 -100
rect 12410 1585 12790 1595
rect 12410 25 12420 1585
rect 12780 25 12790 1585
rect 12410 -725 12790 25
rect 12410 -745 12760 -725
rect 12780 -745 12790 -725
rect 8410 -2375 8420 -815
rect 8780 -2375 8790 -815
rect 8410 -2385 8790 -2375
rect 9210 -815 9590 -805
rect 9210 -2375 9220 -815
rect 9580 -2375 9590 -815
rect 9210 -2385 9590 -2375
rect 10010 -815 10390 -805
rect 10010 -2375 10020 -815
rect 10380 -2375 10390 -815
rect 10010 -2420 10390 -2375
rect 10010 -2500 10020 -2420
rect 10380 -2500 10390 -2420
rect 10010 -2510 10390 -2500
rect 10810 -815 11990 -805
rect 10810 -2375 10820 -815
rect 11180 -2375 11220 -815
rect 11580 -2375 11620 -815
rect 11980 -2375 11990 -815
rect 10810 -2385 11990 -2375
rect 10810 -2420 11190 -2385
rect 10810 -2500 10820 -2420
rect 11180 -2500 11190 -2420
rect 10810 -2510 11190 -2500
rect 11610 -2420 11990 -2385
rect 11610 -2500 11620 -2420
rect 11980 -2500 11990 -2420
rect 11610 -2510 11990 -2500
rect 12410 -815 12790 -745
rect 12410 -2375 12420 -815
rect 12780 -2375 12790 -815
rect 8585 -2625 8625 -2615
rect 8585 -2645 8595 -2625
rect 8615 -2645 8625 -2625
rect 8585 -2670 8625 -2645
rect 8585 -2690 8595 -2670
rect 8615 -2690 8625 -2670
rect 8585 -2700 8625 -2690
rect 7560 -3270 7990 -3260
rect 7560 -3290 7570 -3270
rect 7590 -3290 7990 -3270
rect 7560 -3300 7990 -3290
rect 6810 -4895 6820 -3335
rect 7180 -4895 7190 -3335
rect 6585 -4940 6665 -4930
rect 6585 -4960 6595 -4940
rect 6615 -4960 6635 -4940
rect 6655 -4960 6665 -4940
rect 6585 -4970 6665 -4960
rect 6585 -5125 6625 -5115
rect 6585 -5145 6595 -5125
rect 6615 -5145 6625 -5125
rect 6585 -5170 6625 -5145
rect 6585 -5190 6595 -5170
rect 6615 -5190 6625 -5170
rect 6585 -5200 6625 -5190
rect 6585 -5670 6665 -5660
rect 6585 -5690 6595 -5670
rect 6615 -5690 6635 -5670
rect 6655 -5690 6665 -5670
rect 6585 -5700 6665 -5690
rect 6010 -7295 6020 -5735
rect 6380 -7295 6390 -5735
rect 6010 -7305 6390 -7295
rect 6810 -5735 7190 -4895
rect 6810 -7295 6820 -5735
rect 7180 -7295 7190 -5735
rect 6810 -7305 7190 -7295
rect 7610 -3335 7990 -3325
rect 7610 -4895 7620 -3335
rect 7980 -4895 7990 -3335
rect 7610 -5735 7990 -4895
rect 8410 -3335 8790 -3325
rect 8410 -4895 8420 -3335
rect 8780 -4895 8790 -3335
rect 8410 -4905 8790 -4895
rect 9210 -3335 9590 -3325
rect 9210 -4895 9220 -3335
rect 9580 -4895 9590 -3335
rect 8585 -5125 8625 -5115
rect 8585 -5145 8595 -5125
rect 8615 -5145 8625 -5125
rect 8585 -5170 8625 -5145
rect 8585 -5190 8595 -5170
rect 8615 -5190 8625 -5170
rect 8585 -5200 8625 -5190
rect 7610 -7295 7620 -5735
rect 7980 -7295 7990 -5735
rect 7610 -7305 7990 -7295
rect 8410 -5735 8790 -5725
rect 8410 -7295 8420 -5735
rect 8780 -7295 8790 -5735
rect 8410 -7305 8790 -7295
rect 9210 -5735 9590 -4895
rect 9210 -7295 9220 -5735
rect 9580 -7295 9590 -5735
rect 9210 -7305 9590 -7295
rect 10010 -3335 10390 -3325
rect 10010 -4895 10020 -3335
rect 10380 -4895 10390 -3335
rect 10010 -5645 10390 -4895
rect 10810 -3335 11990 -3325
rect 10810 -4895 10820 -3335
rect 11180 -4895 11220 -3335
rect 11580 -4895 11620 -3335
rect 11980 -4895 11990 -3335
rect 10810 -4905 11990 -4895
rect 10810 -4940 11190 -4905
rect 10810 -5020 10820 -4940
rect 11180 -5020 11190 -4940
rect 10810 -5030 11190 -5020
rect 11610 -4940 11990 -4905
rect 11610 -5020 11620 -4940
rect 11980 -5020 11990 -4940
rect 11610 -5030 11990 -5020
rect 12410 -3335 12790 -2375
rect 13210 1585 13590 1595
rect 13210 25 13220 1585
rect 13580 25 13590 1585
rect 13210 -815 13590 25
rect 14010 1585 14390 1595
rect 14010 25 14020 1585
rect 14380 25 14390 1585
rect 14010 10 14390 25
rect 14810 1585 15190 1595
rect 14810 25 14820 1585
rect 15180 25 15190 1585
rect 14185 -125 14225 -115
rect 14185 -145 14195 -125
rect 14215 -145 14225 -125
rect 14185 -170 14225 -145
rect 14185 -190 14195 -170
rect 14215 -190 14225 -170
rect 14185 -200 14225 -190
rect 13210 -2375 13220 -815
rect 13580 -2375 13590 -815
rect 13210 -2385 13590 -2375
rect 14010 -815 14390 -800
rect 14010 -2375 14020 -815
rect 14380 -2375 14390 -815
rect 14010 -2385 14390 -2375
rect 14810 -815 15190 25
rect 14810 -2375 14820 -815
rect 15180 -2375 15190 -815
rect 14810 -2385 15190 -2375
rect 15610 1585 15990 1595
rect 15610 25 15620 1585
rect 15980 25 15990 1585
rect 15610 -815 15990 25
rect 16410 1585 17190 1595
rect 16410 25 16420 1585
rect 16780 25 16820 1585
rect 17180 25 17190 1585
rect 16410 15 17190 25
rect 18010 1585 18790 1595
rect 18010 25 18020 1585
rect 18380 25 18420 1585
rect 18780 25 18790 1585
rect 18010 15 18790 25
rect 19210 1585 19590 1595
rect 19210 25 19220 1585
rect 19580 25 19590 1585
rect 19210 15 19590 25
rect 20010 1585 20390 1595
rect 20010 25 20020 1585
rect 20380 25 20390 1585
rect 20010 15 20390 25
rect 20810 1585 21190 1595
rect 20810 25 20820 1585
rect 21180 25 21190 1585
rect 20810 15 21190 25
rect 21610 1585 21990 1595
rect 21610 25 21620 1585
rect 21980 25 21990 1585
rect 21610 15 21990 25
rect 22410 1585 22790 1595
rect 22410 25 22420 1585
rect 22780 25 22790 1585
rect 22410 15 22790 25
rect 23210 1585 23990 1595
rect 23210 25 23220 1585
rect 23580 25 23620 1585
rect 23980 25 23990 1585
rect 23210 15 23990 25
rect 16410 -20 16790 15
rect 16410 -100 16420 -20
rect 16780 -100 16790 -20
rect 16410 -110 16790 -100
rect 18410 -20 18790 15
rect 18410 -100 18420 -20
rect 18780 -100 18790 -20
rect 18410 -110 18790 -100
rect 23210 -20 23590 15
rect 23210 -100 23220 -20
rect 23580 -100 23590 -20
rect 23210 -110 23590 -100
rect 20200 -755 21800 -655
rect 20200 -805 20390 -755
rect 21610 -805 21800 -755
rect 15610 -2375 15620 -815
rect 15980 -2375 15990 -815
rect 14185 -2670 14225 -2385
rect 14185 -2690 14195 -2670
rect 14215 -2690 14225 -2670
rect 14185 -2700 14225 -2690
rect 15610 -3220 15990 -2375
rect 16410 -815 17190 -805
rect 16410 -2375 16420 -815
rect 16780 -2375 16820 -815
rect 17180 -2375 17190 -815
rect 16410 -2385 17190 -2375
rect 18010 -815 18790 -805
rect 18010 -2375 18020 -815
rect 18380 -2375 18420 -815
rect 18780 -2375 18790 -815
rect 18010 -2385 18790 -2375
rect 19210 -815 19590 -805
rect 19210 -2375 19220 -815
rect 19580 -2375 19590 -815
rect 19210 -2385 19590 -2375
rect 20010 -815 20390 -805
rect 20010 -2375 20020 -815
rect 20380 -2375 20390 -815
rect 20010 -2385 20390 -2375
rect 20810 -815 21190 -805
rect 20810 -2375 20820 -815
rect 21180 -2375 21190 -815
rect 20810 -2385 21190 -2375
rect 21610 -815 21990 -805
rect 21610 -2375 21620 -815
rect 21980 -2375 21990 -815
rect 21610 -2385 21990 -2375
rect 22410 -815 22790 -805
rect 22410 -2375 22420 -815
rect 22780 -2375 22790 -815
rect 22410 -2385 22790 -2375
rect 23210 -815 23990 -805
rect 23210 -2375 23220 -815
rect 23580 -2375 23620 -815
rect 23980 -2375 23990 -815
rect 23210 -2385 23990 -2375
rect 16410 -2420 16790 -2385
rect 16410 -2500 16420 -2420
rect 16780 -2500 16790 -2420
rect 16410 -2510 16790 -2500
rect 18410 -2420 18790 -2385
rect 18410 -2500 18420 -2420
rect 18780 -2500 18790 -2420
rect 18410 -2510 18790 -2500
rect 23210 -2420 23590 -2385
rect 23210 -2500 23220 -2420
rect 23580 -2500 23590 -2420
rect 23210 -2510 23590 -2500
rect 15610 -3260 17665 -3220
rect 12410 -4895 12420 -3335
rect 12780 -4895 12790 -3335
rect 10585 -5125 10625 -5115
rect 10585 -5145 10595 -5125
rect 10615 -5145 10625 -5125
rect 10585 -5170 10625 -5145
rect 10585 -5190 10595 -5170
rect 10615 -5190 10625 -5170
rect 10585 -5200 10625 -5190
rect 10010 -5665 10020 -5645
rect 10040 -5665 10390 -5645
rect 10010 -5735 10390 -5665
rect 10010 -7295 10020 -5735
rect 10380 -7295 10390 -5735
rect 10010 -7305 10390 -7295
rect 10810 -5735 11990 -5725
rect 10810 -7295 10820 -5735
rect 11180 -7295 11220 -5735
rect 11580 -7295 11620 -5735
rect 11980 -7295 11990 -5735
rect 10810 -7305 11990 -7295
rect 12410 -5735 12790 -4895
rect 12410 -7295 12420 -5735
rect 12780 -7295 12790 -5735
rect 12410 -7305 12790 -7295
rect 13210 -3335 13590 -3325
rect 13210 -4895 13220 -3335
rect 13580 -4895 13590 -3335
rect 13210 -5735 13590 -4895
rect 14010 -3335 14390 -3325
rect 14010 -4895 14020 -3335
rect 14380 -4895 14390 -3335
rect 14010 -4910 14390 -4895
rect 14810 -3335 15190 -3325
rect 14810 -4895 14820 -3335
rect 15180 -4895 15190 -3335
rect 14185 -5125 14225 -5115
rect 14185 -5145 14195 -5125
rect 14215 -5145 14225 -5125
rect 14185 -5170 14225 -5145
rect 14185 -5190 14195 -5170
rect 14215 -5190 14225 -5170
rect 14185 -5200 14225 -5190
rect 13210 -7295 13220 -5735
rect 13580 -7295 13590 -5735
rect 13210 -7305 13590 -7295
rect 14010 -5735 14390 -5720
rect 14010 -7295 14015 -5735
rect 14380 -7295 14390 -5735
rect 14010 -7305 14390 -7295
rect 14810 -5735 15190 -4895
rect 14810 -7295 14820 -5735
rect 15180 -7295 15190 -5735
rect 14810 -7305 15190 -7295
rect 15610 -3335 15990 -3260
rect 20200 -3275 21800 -3175
rect 20200 -3325 20390 -3275
rect 21610 -3325 21800 -3275
rect 15610 -4895 15620 -3335
rect 15980 -4895 15990 -3335
rect 15610 -5735 15990 -4895
rect 16410 -3335 17190 -3325
rect 16410 -4895 16420 -3335
rect 16780 -4895 16820 -3335
rect 17180 -4895 17190 -3335
rect 16410 -4905 17190 -4895
rect 18010 -3335 18790 -3325
rect 18010 -4895 18020 -3335
rect 18380 -4895 18420 -3335
rect 18780 -4895 18790 -3335
rect 18010 -4905 18790 -4895
rect 19210 -3335 19590 -3325
rect 19210 -4895 19220 -3335
rect 19580 -4895 19590 -3335
rect 19210 -4905 19590 -4895
rect 20010 -3335 20390 -3325
rect 20010 -4895 20020 -3335
rect 20380 -4895 20390 -3335
rect 20010 -4905 20390 -4895
rect 20810 -3335 21190 -3325
rect 20810 -4895 20820 -3335
rect 21180 -4895 21190 -3335
rect 20810 -4905 21190 -4895
rect 21610 -3335 21990 -3325
rect 21610 -4895 21620 -3335
rect 21980 -4895 21990 -3335
rect 21610 -4905 21990 -4895
rect 22410 -3335 22790 -3325
rect 22410 -4895 22420 -3335
rect 22780 -4895 22790 -3335
rect 22410 -4905 22790 -4895
rect 23210 -3335 23990 -3325
rect 23210 -4895 23220 -3335
rect 23580 -4895 23620 -3335
rect 23980 -4895 23990 -3335
rect 23210 -4905 23990 -4895
rect 16410 -4940 16790 -4905
rect 16410 -5020 16420 -4940
rect 16780 -5020 16790 -4940
rect 16410 -5030 16790 -5020
rect 18410 -4940 18790 -4905
rect 18410 -5020 18420 -4940
rect 18780 -5020 18790 -4940
rect 18410 -5030 18790 -5020
rect 23210 -4940 23590 -4905
rect 23210 -5020 23220 -4940
rect 23580 -5020 23590 -4940
rect 23210 -5030 23590 -5020
rect 20200 -5675 21800 -5575
rect 20200 -5725 20390 -5675
rect 21610 -5725 21800 -5675
rect 15610 -7295 15620 -5735
rect 15980 -7295 15990 -5735
rect 15610 -7305 15990 -7295
rect 16410 -5735 17190 -5725
rect 16410 -7295 16420 -5735
rect 16780 -7295 16820 -5735
rect 17180 -7295 17190 -5735
rect 16410 -7305 17190 -7295
rect 18010 -5735 18790 -5725
rect 18010 -7295 18020 -5735
rect 18380 -7295 18420 -5735
rect 18780 -7295 18790 -5735
rect 18010 -7305 18790 -7295
rect 19210 -5735 19590 -5725
rect 19210 -7295 19220 -5735
rect 19580 -7295 19590 -5735
rect 19210 -7305 19590 -7295
rect 20010 -5735 20390 -5725
rect 20010 -7295 20020 -5735
rect 20380 -7295 20390 -5735
rect 20010 -7305 20390 -7295
rect 20810 -5735 21190 -5725
rect 20810 -7295 20820 -5735
rect 21180 -7295 21190 -5735
rect 20810 -7305 21190 -7295
rect 21610 -5735 21990 -5725
rect 21610 -7295 21620 -5735
rect 21980 -7295 21990 -5735
rect 21610 -7305 21990 -7295
rect 22410 -5735 22790 -5725
rect 22410 -7295 22420 -5735
rect 22780 -7295 22790 -5735
rect 22410 -7305 22790 -7295
rect 23210 -5735 23990 -5725
rect 23210 -7295 23220 -5735
rect 23580 -7295 23620 -5735
rect 23980 -7295 23990 -5735
rect 23210 -7305 23990 -7295
rect -390 -7340 -10 -7305
rect -390 -7420 -380 -7340
rect -20 -7420 -10 -7340
rect 2180 -7330 2220 -7325
rect 2180 -7350 2190 -7330
rect 2210 -7350 2220 -7330
rect 2180 -7370 2220 -7350
rect 2180 -7390 2190 -7370
rect 2210 -7390 2220 -7370
rect 4580 -7360 4620 -7305
rect 4580 -7380 4590 -7360
rect 4610 -7380 4620 -7360
rect 4580 -7390 4620 -7380
rect 6180 -7330 6220 -7325
rect 6180 -7350 6190 -7330
rect 6210 -7350 6220 -7330
rect 6180 -7370 6220 -7350
rect 6180 -7390 6190 -7370
rect 6210 -7390 6220 -7370
rect 2180 -7400 2220 -7390
rect 6180 -7400 6220 -7390
rect 7200 -7340 7600 -7330
rect -390 -7430 -10 -7420
rect 7200 -7420 7210 -7340
rect 7590 -7420 7600 -7340
rect 7200 -7455 7600 -7420
rect 8000 -7340 8400 -7330
rect 8000 -7420 8010 -7340
rect 8390 -7420 8400 -7340
rect 8580 -7360 8620 -7305
rect 8580 -7380 8590 -7360
rect 8610 -7380 8620 -7360
rect 8580 -7390 8620 -7380
rect 8800 -7340 9200 -7330
rect 8000 -7455 8400 -7420
rect 8800 -7420 8810 -7340
rect 9190 -7420 9200 -7340
rect 8800 -7455 9200 -7420
rect 9600 -7340 10000 -7330
rect 9600 -7420 9610 -7340
rect 9990 -7420 10000 -7340
rect 9600 -7455 10000 -7420
rect 10810 -7340 11190 -7305
rect 10810 -7420 10820 -7340
rect 11180 -7420 11190 -7340
rect 10810 -7430 11190 -7420
rect 11610 -7340 11990 -7305
rect 11610 -7420 11620 -7340
rect 11980 -7420 11990 -7340
rect 11610 -7430 11990 -7420
rect 12800 -7340 13200 -7330
rect 12800 -7420 12810 -7340
rect 13190 -7420 13200 -7340
rect 12800 -7455 13200 -7420
rect 13600 -7340 14000 -7330
rect 13600 -7420 13610 -7340
rect 13990 -7420 14000 -7340
rect 14185 -7360 14225 -7305
rect 14185 -7380 14195 -7360
rect 14215 -7380 14225 -7360
rect 14185 -7390 14225 -7380
rect 16410 -7340 16790 -7305
rect 13600 -7455 14000 -7420
rect 16410 -7420 16420 -7340
rect 16780 -7420 16790 -7340
rect 16410 -7430 16790 -7420
rect 18410 -7340 18790 -7305
rect 18410 -7420 18420 -7340
rect 18780 -7420 18790 -7340
rect 18410 -7430 18790 -7420
rect 19600 -7340 20000 -7330
rect 19600 -7420 19610 -7340
rect 19990 -7420 20000 -7340
rect 19600 -7455 20000 -7420
rect 20400 -7340 20800 -7330
rect 20400 -7420 20410 -7340
rect 20790 -7420 20800 -7340
rect 20400 -7455 20800 -7420
rect 21200 -7340 21600 -7330
rect 21200 -7420 21210 -7340
rect 21590 -7420 21600 -7340
rect 21200 -7455 21600 -7420
rect 22000 -7340 22400 -7330
rect 22000 -7420 22010 -7340
rect 22390 -7420 22400 -7340
rect 22000 -7455 22400 -7420
rect 23210 -7340 23590 -7305
rect 23210 -7420 23220 -7340
rect 23580 -7420 23590 -7340
rect 23210 -7430 23590 -7420
rect 7200 -7555 22400 -7455
<< viali >>
rect 5385 2040 5405 2060
rect 14195 1855 14215 1875
rect 1390 1785 1410 1805
rect 3210 1730 3590 1820
rect 3780 1785 3800 1805
rect 8190 1790 8210 1810
rect -780 25 -420 1585
rect -380 25 -20 1585
rect 1220 25 1580 1585
rect 1390 -215 1410 -195
rect -780 -2375 -420 -815
rect -380 -2375 -20 -815
rect 1220 -2375 1580 -815
rect 3780 -215 3800 -195
rect 3210 -670 3590 -575
rect 2190 -2645 2210 -2625
rect -780 -4895 -420 -3335
rect -380 -4895 -20 -3335
rect 5220 25 5580 1585
rect 5960 -80 5980 -60
rect 5385 -210 5405 -190
rect 5960 -730 5980 -710
rect 5220 -2375 5580 -815
rect 6420 -80 6440 -60
rect 6420 -730 6440 -710
rect 7220 -670 7580 -575
rect 4575 -2645 4595 -2625
rect 6595 -2645 6615 -2625
rect 6020 -3265 6380 -3185
rect 4420 -4895 4780 -3335
rect -780 -7295 -420 -5735
rect -380 -7295 -20 -5735
rect 2190 -5145 2210 -5125
rect 4575 -5145 4595 -5125
rect 4420 -7295 4780 -5735
rect 8190 -210 8210 -190
rect 9220 25 9580 1585
rect 10020 25 10380 1585
rect 10820 25 11180 1585
rect 11220 25 11580 1585
rect 11620 25 11980 1585
rect 9220 -2375 9580 -815
rect 10020 -2375 10380 -815
rect 10820 -2375 11180 -815
rect 11220 -2375 11580 -815
rect 11620 -2375 11980 -815
rect 8595 -2645 8615 -2625
rect 6635 -4960 6655 -4940
rect 6595 -5145 6615 -5125
rect 6635 -5690 6655 -5670
rect 8420 -4895 8780 -3335
rect 8595 -5145 8615 -5125
rect 8420 -7295 8780 -5735
rect 10820 -4895 11180 -3335
rect 11220 -4895 11580 -3335
rect 11620 -4895 11980 -3335
rect 14020 25 14380 1585
rect 14195 -145 14215 -125
rect 14020 -2375 14380 -815
rect 16420 25 16780 1585
rect 16820 25 17180 1585
rect 20820 25 21180 1585
rect 16420 -2375 16780 -815
rect 16820 -2375 17180 -815
rect 20820 -2375 21180 -815
rect 10595 -5145 10615 -5125
rect 10820 -7295 11180 -5735
rect 11220 -7295 11580 -5735
rect 11620 -7295 11980 -5735
rect 14020 -4895 14380 -3335
rect 14195 -5145 14215 -5125
rect 14015 -7295 14380 -5735
rect 16420 -4895 16780 -3335
rect 16820 -4895 17180 -3335
rect 20820 -4895 21180 -3335
rect 16420 -7295 16780 -5735
rect 16820 -7295 17180 -5735
rect 20820 -7295 21180 -5735
rect 2190 -7350 2210 -7330
rect 6190 -7350 6210 -7330
<< metal1 >>
rect -800 2060 24000 2595
rect -800 2040 5385 2060
rect 5405 2040 24000 2060
rect -800 1875 24000 2040
rect -800 1855 14195 1875
rect 14215 1855 24000 1875
rect -800 1820 24000 1855
rect -800 1805 3210 1820
rect -800 1785 1390 1805
rect 1410 1785 3210 1805
rect -800 1730 3210 1785
rect 3590 1810 24000 1820
rect 3590 1805 8190 1810
rect 3590 1785 3780 1805
rect 3800 1790 8190 1805
rect 8210 1790 24000 1810
rect 3800 1785 24000 1790
rect 3590 1730 24000 1785
rect -800 1595 24000 1730
rect -800 1585 5785 1595
rect -800 25 -780 1585
rect -420 25 -380 1585
rect -20 25 1220 1585
rect 1580 25 5220 1585
rect 5580 25 5785 1585
rect -800 -190 5785 25
rect 6610 1585 24000 1595
rect 6610 25 9220 1585
rect 9580 25 10020 1585
rect 10380 25 10820 1585
rect 11180 25 11220 1585
rect 11580 25 11620 1585
rect 11980 25 14020 1585
rect 14380 25 16420 1585
rect 16780 25 16820 1585
rect 17180 25 20820 1585
rect 21180 25 24000 1585
rect -800 -195 5385 -190
rect -800 -215 1390 -195
rect 1410 -215 3780 -195
rect 3800 -210 5385 -195
rect 5405 -210 5785 -190
rect 3800 -215 5785 -210
rect -800 -575 5785 -215
rect -800 -670 3210 -575
rect 3590 -670 5785 -575
rect -800 -815 5785 -670
rect 5930 -60 6470 5
rect 5930 -80 5960 -60
rect 5980 -80 6420 -60
rect 6440 -80 6470 -60
rect 5930 -710 6470 -80
rect 5930 -730 5960 -710
rect 5980 -730 6420 -710
rect 6440 -730 6470 -710
rect 5930 -780 6470 -730
rect 6610 -125 24000 25
rect 6610 -145 14195 -125
rect 14215 -145 24000 -125
rect 6610 -190 24000 -145
rect 6610 -210 8190 -190
rect 8210 -210 24000 -190
rect 6610 -575 24000 -210
rect 6610 -670 7220 -575
rect 7580 -670 24000 -575
rect -800 -2375 -780 -815
rect -420 -2375 -380 -815
rect -20 -2375 1220 -815
rect 1580 -2375 5220 -815
rect 5580 -2375 5785 -815
rect -800 -2385 5785 -2375
rect 2010 -2625 2390 -2615
rect 2010 -2645 2190 -2625
rect 2210 -2645 2390 -2625
rect 2010 -3325 2390 -2645
rect 4410 -2625 4790 -2615
rect 4410 -2645 4575 -2625
rect 4595 -2645 4790 -2625
rect 4410 -3325 4790 -2645
rect 6010 -3185 6390 -780
rect 6610 -815 24000 -670
rect 6610 -2375 9220 -815
rect 9580 -2375 10020 -815
rect 10380 -2375 10820 -815
rect 11180 -2375 11220 -815
rect 11580 -2375 11620 -815
rect 11980 -2375 14020 -815
rect 14380 -2375 16420 -815
rect 16780 -2375 16820 -815
rect 17180 -2375 20820 -815
rect 21180 -2375 24000 -815
rect 6610 -2385 24000 -2375
rect 6010 -3265 6020 -3185
rect 6380 -3265 6390 -3185
rect 6010 -3275 6390 -3265
rect 6420 -2625 6780 -2615
rect 6420 -2645 6595 -2625
rect 6615 -2645 6780 -2625
rect 6420 -3325 6780 -2645
rect 8410 -2625 8790 -2615
rect 8410 -2645 8595 -2625
rect 8615 -2645 8790 -2625
rect 8410 -3325 8790 -2645
rect 12410 -3325 12790 -2385
rect 14180 -2705 14230 -2655
rect 15610 -3220 15990 -2385
rect 15610 -3260 17665 -3220
rect 15610 -3325 15990 -3260
rect 20800 -3325 21200 -2385
rect -800 -3335 24000 -3325
rect -800 -4895 -780 -3335
rect -420 -4895 -380 -3335
rect -20 -4895 4420 -3335
rect 4780 -4895 8420 -3335
rect 8780 -4895 10820 -3335
rect 11180 -4895 11220 -3335
rect 11580 -4895 11620 -3335
rect 11980 -4895 14020 -3335
rect 14380 -4895 16420 -3335
rect 16780 -4895 16820 -3335
rect 17180 -4895 20820 -3335
rect 21180 -4895 24000 -3335
rect -800 -4940 24000 -4895
rect -800 -4960 6635 -4940
rect 6655 -4960 24000 -4940
rect -800 -5125 24000 -4960
rect -800 -5145 2190 -5125
rect 2210 -5145 4575 -5125
rect 4595 -5145 6595 -5125
rect 6615 -5145 8595 -5125
rect 8615 -5145 10595 -5125
rect 10615 -5145 14195 -5125
rect 14215 -5145 24000 -5125
rect -800 -5670 24000 -5145
rect -800 -5690 6635 -5670
rect 6655 -5690 24000 -5670
rect -800 -5735 24000 -5690
rect -800 -7295 -780 -5735
rect -420 -7295 -380 -5735
rect -20 -7295 4420 -5735
rect 4780 -7295 8420 -5735
rect 8780 -7295 10820 -5735
rect 11180 -7295 11220 -5735
rect 11580 -7295 11620 -5735
rect 11980 -7295 14015 -5735
rect 14380 -7295 16420 -5735
rect 16780 -7295 16820 -5735
rect 17180 -7295 20820 -5735
rect 21180 -7295 24000 -5735
rect -800 -7305 24000 -7295
rect 2010 -7330 2390 -7305
rect 2010 -7350 2190 -7330
rect 2210 -7350 2390 -7330
rect 2010 -7415 2390 -7350
rect 6010 -7330 6390 -7305
rect 10000 -7310 10430 -7305
rect 20800 -7315 21200 -7305
rect 6010 -7350 6190 -7330
rect 6210 -7350 6390 -7330
rect 6010 -7415 6390 -7350
<< end >>
