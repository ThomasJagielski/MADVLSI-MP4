magic
tech sky130A
timestamp 1617421225
<< nwell >>
rect -615 -160 15825 1710
<< pmos >>
rect 205 0 605 1600
rect 1005 0 1405 1600
rect 1805 0 2205 1600
rect 2605 0 3005 1600
rect 3405 0 3805 1600
rect 4205 0 4605 1600
rect 5005 0 5405 1600
rect 5805 0 6205 1600
rect 6605 0 7005 1600
rect 7405 0 7805 1600
rect 8205 0 8605 1600
rect 9005 0 9405 1600
rect 9805 0 10205 1600
rect 10605 0 11005 1600
rect 11405 0 11805 1600
rect 12205 0 12605 1600
rect 13005 0 13405 1600
rect 13805 0 14205 1600
rect 14605 0 15005 1600
<< pdiff >>
rect -195 1585 205 1600
rect -195 15 -180 1585
rect 190 15 205 1585
rect -195 0 205 15
rect 605 1585 1005 1600
rect 605 15 620 1585
rect 990 15 1005 1585
rect 605 0 1005 15
rect 1405 1585 1805 1600
rect 1405 15 1420 1585
rect 1790 15 1805 1585
rect 1405 0 1805 15
rect 2205 1585 2605 1600
rect 2205 15 2220 1585
rect 2590 15 2605 1585
rect 2205 0 2605 15
rect 3005 1585 3405 1600
rect 3005 15 3020 1585
rect 3395 15 3405 1585
rect 3005 0 3405 15
rect 3805 1585 4205 1600
rect 3805 15 3820 1585
rect 4190 15 4205 1585
rect 3805 0 4205 15
rect 4605 1585 5005 1600
rect 4605 15 4620 1585
rect 4990 15 5005 1585
rect 4605 0 5005 15
rect 5405 1585 5805 1600
rect 5405 15 5420 1585
rect 5790 15 5805 1585
rect 5405 0 5805 15
rect 6205 1585 6605 1600
rect 6205 15 6220 1585
rect 6590 15 6605 1585
rect 6205 0 6605 15
rect 7005 1585 7405 1600
rect 7005 15 7020 1585
rect 7390 15 7405 1585
rect 7005 0 7405 15
rect 7805 1585 8205 1600
rect 7805 15 7820 1585
rect 8190 15 8205 1585
rect 7805 0 8205 15
rect 8605 1585 9005 1600
rect 8605 15 8620 1585
rect 8990 15 9005 1585
rect 8605 0 9005 15
rect 9405 1585 9805 1600
rect 9405 15 9420 1585
rect 9790 15 9805 1585
rect 9405 0 9805 15
rect 10205 1585 10605 1600
rect 10205 15 10220 1585
rect 10590 15 10605 1585
rect 10205 0 10605 15
rect 11005 1585 11405 1600
rect 11005 15 11020 1585
rect 11390 15 11405 1585
rect 11005 0 11405 15
rect 11805 1585 12205 1600
rect 11805 15 11820 1585
rect 12190 15 12205 1585
rect 11805 0 12205 15
rect 12605 1585 13005 1600
rect 12605 15 12620 1585
rect 12990 15 13005 1585
rect 12605 0 13005 15
rect 13405 1585 13805 1600
rect 13405 15 13420 1585
rect 13790 15 13805 1585
rect 13405 0 13805 15
rect 14205 1585 14605 1600
rect 14205 15 14220 1585
rect 14590 15 14605 1585
rect 14205 0 14605 15
rect 15005 1585 15405 1600
rect 15005 15 15020 1585
rect 15390 15 15405 1585
rect 15005 0 15405 15
<< pdiffc >>
rect -180 15 190 1585
rect 620 15 990 1585
rect 1420 15 1790 1585
rect 2220 15 2590 1585
rect 3020 15 3395 1585
rect 3820 15 4190 1585
rect 4620 15 4990 1585
rect 5420 15 5790 1585
rect 6220 15 6590 1585
rect 7020 15 7390 1585
rect 7820 15 8190 1585
rect 8620 15 8990 1585
rect 9420 15 9790 1585
rect 10220 15 10590 1585
rect 11020 15 11390 1585
rect 11820 15 12190 1585
rect 12620 15 12990 1585
rect 13420 15 13790 1585
rect 14220 15 14590 1585
rect 15020 15 15390 1585
<< nsubdiff >>
rect 1560 1675 1610 1690
rect 1560 1655 1575 1675
rect 1595 1655 1610 1675
rect 3575 1665 3625 1680
rect 1560 1640 1610 1655
rect 3575 1645 3590 1665
rect 3610 1645 3625 1665
rect 6350 1665 6400 1680
rect 3575 1630 3625 1645
rect 6350 1645 6365 1665
rect 6385 1645 6400 1665
rect 6350 1630 6400 1645
rect 7960 1665 8010 1680
rect 7960 1645 7975 1665
rect 7995 1645 8010 1665
rect 7960 1630 8010 1645
rect 9580 1665 9630 1680
rect 9580 1645 9595 1665
rect 9615 1645 9630 1665
rect 12390 1665 12440 1680
rect 9580 1630 9630 1645
rect 12390 1645 12405 1665
rect 12425 1645 12440 1665
rect 12390 1630 12440 1645
rect -595 1585 -195 1600
rect -595 15 -580 1585
rect -210 15 -195 1585
rect -595 0 -195 15
rect 15405 1585 15805 1600
rect 15405 15 15420 1585
rect 15790 15 15805 1585
rect 15405 0 15805 15
rect 2775 -85 2825 -70
rect 2775 -105 2790 -85
rect 2810 -105 2825 -85
rect 2775 -120 2825 -105
rect 3575 -85 3625 -70
rect 3575 -105 3590 -85
rect 3610 -105 3625 -85
rect 3575 -120 3625 -105
rect 6375 -60 6425 -45
rect 6375 -80 6390 -60
rect 6410 -80 6425 -60
rect 6375 -95 6425 -80
rect 7550 -60 7600 -45
rect 9585 -60 9635 -45
rect 7550 -80 7565 -60
rect 7585 -80 7600 -60
rect 7550 -95 7600 -80
rect 9585 -80 9600 -60
rect 9620 -80 9635 -60
rect 9585 -95 9635 -80
rect 12380 -85 12430 -70
rect 12380 -105 12395 -85
rect 12415 -105 12430 -85
rect 12380 -120 12430 -105
<< nsubdiffcont >>
rect 1575 1655 1595 1675
rect 3590 1645 3610 1665
rect 6365 1645 6385 1665
rect 7975 1645 7995 1665
rect 9595 1645 9615 1665
rect 12405 1645 12425 1665
rect -580 15 -210 1585
rect 15420 15 15790 1585
rect 2790 -105 2810 -85
rect 3590 -105 3610 -85
rect 6390 -80 6410 -60
rect 7565 -80 7585 -60
rect 9600 -80 9620 -60
rect 12395 -105 12415 -85
<< poly >>
rect 35 1645 75 1655
rect 35 1630 45 1645
rect -190 1625 45 1630
rect 65 1630 75 1645
rect 835 1645 875 1655
rect 835 1630 845 1645
rect 65 1625 845 1630
rect 865 1630 875 1645
rect 1635 1645 1675 1655
rect 1635 1630 1645 1645
rect 865 1625 1645 1630
rect 1665 1630 1675 1645
rect 2435 1645 2475 1655
rect 2435 1630 2445 1645
rect 1665 1625 2445 1630
rect 2465 1630 2475 1645
rect 4435 1645 4475 1655
rect 2465 1625 3005 1630
rect -190 1615 3005 1625
rect 4435 1625 4445 1645
rect 4465 1625 4475 1645
rect 11635 1645 11675 1655
rect 4435 1615 4475 1625
rect 11635 1625 11645 1645
rect 11665 1625 11675 1645
rect 13625 1645 13665 1655
rect 13625 1630 13635 1645
rect 11635 1615 11675 1625
rect 13005 1625 13635 1630
rect 13655 1630 13665 1645
rect 14425 1645 14465 1655
rect 14425 1630 14435 1645
rect 13655 1625 14435 1630
rect 14455 1630 14465 1645
rect 15235 1645 15275 1655
rect 15235 1630 15245 1645
rect 14455 1625 15245 1630
rect 15265 1630 15275 1645
rect 15265 1625 15400 1630
rect 13005 1615 15400 1625
rect 205 1600 605 1615
rect 1005 1600 1405 1615
rect 1805 1600 2205 1615
rect 2605 1600 3005 1615
rect 3405 1600 3805 1615
rect 4205 1600 4605 1615
rect 5005 1600 5405 1615
rect 5805 1600 6205 1615
rect 6605 1600 7005 1615
rect 7405 1600 7805 1615
rect 8205 1600 8605 1615
rect 9005 1600 9405 1615
rect 9805 1600 10205 1615
rect 10605 1600 11005 1615
rect 11405 1600 11805 1615
rect 12205 1600 12605 1615
rect 13005 1600 13405 1615
rect 13805 1600 14205 1615
rect 14605 1600 15005 1615
rect 205 -15 605 0
rect 1005 -15 1405 0
rect 1805 -15 2205 0
rect 2605 -15 3005 0
rect 3405 -45 3805 0
rect 4205 -15 4605 0
rect 5005 -45 5405 0
rect 5805 -20 6205 0
rect 6605 -20 7005 0
rect 7405 -20 7805 0
rect 8205 -20 8605 0
rect 9005 -20 9405 0
rect 9805 -20 10205 0
rect 5805 -35 10205 -20
rect 10605 -45 11005 0
rect 11405 -15 11805 0
rect 12205 -45 12605 0
rect 13005 -15 13405 0
rect 13805 -15 14205 0
rect 14605 -15 15005 0
rect 3405 -55 5405 -45
rect 3405 -60 4970 -55
rect 4960 -75 4970 -60
rect 4990 -60 5405 -55
rect 4990 -75 5000 -60
rect 4960 -85 5000 -75
rect 4960 -175 4975 -85
rect 10605 -55 12605 -45
rect 10605 -60 11020 -55
rect 8035 -70 8075 -60
rect 8035 -90 8045 -70
rect 8065 -90 8075 -70
rect 8035 -100 8075 -90
rect 11010 -75 11020 -60
rect 11040 -60 12605 -55
rect 11040 -75 11050 -60
rect 11010 -85 11050 -75
rect 4960 -185 5000 -175
rect 4960 -205 4970 -185
rect 4990 -205 5000 -185
rect 4960 -215 5000 -205
rect 8035 -235 8050 -100
rect 8035 -245 8075 -235
rect 8035 -265 8045 -245
rect 8065 -265 8075 -245
rect 8035 -275 8075 -265
<< polycont >>
rect 45 1625 65 1645
rect 845 1625 865 1645
rect 1645 1625 1665 1645
rect 2445 1625 2465 1645
rect 4445 1625 4465 1645
rect 11645 1625 11665 1645
rect 13635 1625 13655 1645
rect 14435 1625 14455 1645
rect 15245 1625 15265 1645
rect 4970 -75 4990 -55
rect 8045 -90 8065 -70
rect 11020 -75 11040 -55
rect 4970 -205 4990 -185
rect 8045 -265 8065 -245
<< locali >>
rect 3010 1765 13000 1785
rect 1565 1675 1605 1685
rect 1565 1655 1575 1675
rect 1595 1655 1605 1675
rect 35 1645 75 1655
rect 35 1625 45 1645
rect 65 1625 75 1645
rect 35 1615 75 1625
rect 835 1645 875 1655
rect 835 1625 845 1645
rect 865 1625 875 1645
rect 835 1615 875 1625
rect 1565 1615 1605 1655
rect 1635 1645 1675 1655
rect 1635 1625 1645 1645
rect 1665 1625 1675 1645
rect 1635 1615 1675 1625
rect 2435 1645 2475 1655
rect 2435 1625 2445 1645
rect 2465 1625 2475 1645
rect 2435 1615 2475 1625
rect -190 1595 200 1615
rect -590 1585 200 1595
rect -590 15 -580 1585
rect -210 15 -180 1585
rect 190 15 200 1585
rect -590 5 200 15
rect 610 1585 1000 1615
rect 610 15 620 1585
rect 990 15 1000 1585
rect 610 5 1000 15
rect 1410 1585 1800 1615
rect 1410 15 1420 1585
rect 1790 15 1800 1585
rect 1410 0 1800 15
rect 2210 1585 2600 1615
rect 2210 15 2220 1585
rect 2590 15 2600 1585
rect 2210 5 2600 15
rect 3010 1585 3400 1765
rect 3810 1740 12195 1745
rect 3810 1725 12200 1740
rect 3580 1665 3620 1675
rect 3580 1645 3590 1665
rect 3610 1645 3620 1665
rect 3580 1635 3620 1645
rect 3010 15 3020 1585
rect 3395 15 3400 1585
rect 3010 -30 3400 15
rect 3810 1585 4200 1725
rect 4435 1685 4475 1695
rect 4435 1665 4445 1685
rect 4465 1665 4475 1685
rect 4435 1645 4475 1665
rect 4435 1625 4445 1645
rect 4465 1625 4475 1645
rect 4435 1615 4475 1625
rect 6355 1665 6395 1675
rect 6355 1645 6365 1665
rect 6385 1645 6395 1665
rect 6355 1595 6395 1645
rect 3810 15 3820 1585
rect 4190 15 4200 1585
rect 3810 0 4200 15
rect 4610 1585 5000 1595
rect 4610 15 4620 1585
rect 4990 15 5000 1585
rect -615 -50 3400 -30
rect 4610 -45 5000 15
rect 4960 -55 5000 -45
rect 4960 -75 4970 -55
rect 4990 -75 5000 -55
rect 2780 -85 2820 -75
rect 2780 -105 2790 -85
rect 2810 -105 2820 -85
rect 2780 -115 2820 -105
rect 3580 -85 3620 -75
rect 4960 -85 5000 -75
rect 5410 1585 5800 1595
rect 5410 15 5420 1585
rect 5790 15 5800 1585
rect 3580 -105 3590 -85
rect 3610 -105 3620 -85
rect 3580 -115 3620 -105
rect 5410 -135 5800 15
rect 6210 1585 6600 1595
rect 6210 15 6220 1585
rect 6590 15 6600 1585
rect 6210 5 6600 15
rect 7010 1585 7400 1725
rect 7965 1665 8005 1675
rect 7965 1645 7975 1665
rect 7995 1645 8005 1665
rect 7965 1635 8005 1645
rect 7010 15 7020 1585
rect 7390 15 7400 1585
rect 6380 -60 6420 5
rect 7010 0 7400 15
rect 7810 1585 8200 1595
rect 7810 15 7820 1585
rect 8190 15 8200 1585
rect 6380 -80 6390 -60
rect 6410 -80 6420 -60
rect 6380 -90 6420 -80
rect 7555 -60 7595 -50
rect 7810 -60 8200 15
rect 8610 1585 9000 1725
rect 11635 1685 11675 1695
rect 9585 1665 9625 1675
rect 9585 1645 9595 1665
rect 9615 1645 9625 1665
rect 9585 1595 9625 1645
rect 11635 1665 11645 1685
rect 11665 1665 11675 1685
rect 11635 1645 11675 1665
rect 11635 1625 11645 1645
rect 11665 1625 11675 1645
rect 11635 1615 11675 1625
rect 8610 15 8620 1585
rect 8990 15 9000 1585
rect 8610 0 9000 15
rect 9410 1585 9800 1595
rect 9410 15 9420 1585
rect 9790 15 9800 1585
rect 9410 5 9800 15
rect 10210 1585 10600 1595
rect 10210 15 10220 1585
rect 10590 15 10600 1585
rect 9590 -60 9630 5
rect 7555 -80 7565 -60
rect 7585 -80 7595 -60
rect 7555 -90 7595 -80
rect 8035 -70 8075 -60
rect 8035 -90 8045 -70
rect 8065 -90 8075 -70
rect 9590 -80 9600 -60
rect 9620 -80 9630 -60
rect 9590 -90 9630 -80
rect 8035 -100 8075 -90
rect -615 -145 5800 -135
rect 10210 -145 10600 15
rect -615 -155 10600 -145
rect 5410 -165 10600 -155
rect 11010 1585 11400 1595
rect 11010 15 11020 1585
rect 11390 15 11400 1585
rect 11010 -45 11400 15
rect 11810 1585 12200 1725
rect 12395 1665 12435 1675
rect 12395 1645 12405 1665
rect 12425 1645 12435 1665
rect 12395 1635 12435 1645
rect 11810 15 11820 1585
rect 12190 15 12200 1585
rect 11810 5 12200 15
rect 12610 1585 13000 1765
rect 13625 1645 13665 1655
rect 13625 1625 13635 1645
rect 13655 1625 13665 1645
rect 13625 1615 13665 1625
rect 14425 1645 14465 1655
rect 14425 1625 14435 1645
rect 14455 1625 14465 1645
rect 14425 1615 14465 1625
rect 15235 1645 15275 1655
rect 15235 1625 15245 1645
rect 15265 1625 15275 1645
rect 15235 1615 15275 1625
rect 12610 15 12620 1585
rect 12990 15 13000 1585
rect 12610 5 13000 15
rect 13410 1585 13800 1595
rect 13410 15 13420 1585
rect 13790 15 13800 1585
rect 13410 0 13800 15
rect 14210 1585 14600 1615
rect 14210 15 14220 1585
rect 14590 15 14600 1585
rect 14210 5 14600 15
rect 15010 1595 15400 1615
rect 15010 1585 15800 1595
rect 15010 15 15020 1585
rect 15390 15 15420 1585
rect 15790 15 15800 1585
rect 15010 5 15800 15
rect 11010 -55 11050 -45
rect 11010 -75 11020 -55
rect 11040 -75 11050 -55
rect 11010 -85 11050 -75
rect 12385 -85 12425 -75
rect 4960 -185 5000 -175
rect 4960 -195 4970 -185
rect -615 -205 4970 -195
rect 4990 -195 5000 -185
rect 11010 -195 11030 -85
rect 12385 -105 12395 -85
rect 12415 -105 12425 -85
rect 12385 -115 12425 -105
rect 4990 -205 11030 -195
rect -615 -215 11030 -205
rect -615 -245 8075 -235
rect -615 -255 8045 -245
rect 8035 -265 8045 -255
rect 8065 -265 8075 -245
rect 8035 -275 8075 -265
<< viali >>
rect -580 15 -210 1585
rect -180 15 190 1585
rect 620 15 990 1585
rect 1420 15 1790 1585
rect 2220 15 2590 1585
rect 3590 1645 3610 1665
rect 4445 1665 4465 1685
rect 2790 -105 2810 -85
rect 3590 -105 3610 -85
rect 6220 15 6590 1585
rect 7975 1645 7995 1665
rect 11645 1665 11665 1685
rect 9420 15 9790 1585
rect 7565 -80 7585 -60
rect 12405 1645 12425 1665
rect 13420 15 13790 1585
rect 14220 15 14590 1585
rect 15020 15 15390 1585
rect 15420 15 15790 1585
rect 12395 -105 12415 -85
<< metal1 >>
rect 4435 1685 4475 1695
rect 3580 1665 3620 1675
rect 3580 1645 3590 1665
rect 3610 1645 3620 1665
rect 3580 1595 3620 1645
rect 4435 1665 4445 1685
rect 4465 1665 4475 1685
rect 11635 1685 11675 1695
rect 4435 1595 4475 1665
rect 7965 1665 8005 1675
rect 7965 1645 7975 1665
rect 7995 1645 8005 1665
rect 7965 1595 8005 1645
rect 11635 1665 11645 1685
rect 11665 1665 11675 1685
rect 11635 1595 11675 1665
rect 12395 1665 12435 1675
rect 12395 1645 12405 1665
rect 12425 1645 12435 1665
rect 12395 1595 12435 1645
rect -595 1585 15805 1595
rect -595 15 -580 1585
rect -210 15 -180 1585
rect 190 15 620 1585
rect 990 15 1420 1585
rect 1790 15 2220 1585
rect 2590 15 6220 1585
rect 6590 15 9420 1585
rect 9790 15 13420 1585
rect 13790 15 14220 1585
rect 14590 15 15020 1585
rect 15390 15 15420 1585
rect 15790 15 15805 1585
rect -595 5 15805 15
rect 2780 -85 2820 5
rect 2780 -105 2790 -85
rect 2810 -105 2820 -85
rect 2780 -115 2820 -105
rect 3580 -85 3620 5
rect 3580 -105 3590 -85
rect 3610 -105 3620 -85
rect 7555 -60 7595 5
rect 7555 -80 7565 -60
rect 7585 -80 7595 -60
rect 7555 -90 7595 -80
rect 12385 -85 12425 5
rect 3580 -115 3620 -105
rect 12385 -105 12395 -85
rect 12415 -105 12425 -85
rect 12385 -115 12425 -105
<< labels >>
rlabel metal1 -595 800 -595 800 7 VP
rlabel locali -615 -40 -615 -40 7 Vout
rlabel locali -615 -145 -615 -145 7 Iin
<< end >>
