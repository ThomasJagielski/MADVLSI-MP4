magic
tech sky130A
timestamp 1617545523
<< nmos >>
rect -1900 0 -1500 1600
rect -1200 0 -800 1600
rect -500 0 -100 1600
rect 200 0 600 1600
rect 900 0 1300 1600
rect 1600 0 2000 1600
rect 2300 0 2700 1600
rect 3000 0 3400 1600
rect 3700 0 4100 1600
rect 4400 0 4800 1600
rect 5100 0 5500 1600
rect 5800 0 6200 1600
rect 6500 0 6900 1600
rect 7200 0 7600 1600
rect 7900 0 8300 1600
rect 8600 0 9000 1600
rect 9300 0 9700 1600
rect 10000 0 10400 1600
rect 10700 0 11100 1600
rect -1900 -2000 -1500 -400
rect -1200 -2000 -800 -400
rect -500 -2000 -100 -400
rect 200 -2000 600 -400
rect 900 -2000 1300 -400
rect 1600 -2000 2000 -400
rect 2300 -2000 2700 -400
rect 3000 -2000 3400 -400
rect 3700 -2000 4100 -400
rect 4400 -2000 4800 -400
rect 5100 -2000 5500 -400
rect 5800 -2000 6200 -400
rect 6500 -2000 6900 -400
rect 7200 -2000 7600 -400
rect 7900 -2000 8300 -400
rect 8600 -2000 9000 -400
rect 9300 -2000 9700 -400
rect 10000 -2000 10400 -400
rect 10700 -2000 11100 -400
rect -1900 -4000 -1500 -2400
rect -1200 -4000 -800 -2400
rect -500 -4000 -100 -2400
rect 200 -4000 600 -2400
rect 900 -4000 1300 -2400
rect 1600 -4000 2000 -2400
rect 2300 -4000 2700 -2400
rect 3000 -4000 3400 -2400
rect 3700 -4000 4100 -2400
rect 4400 -4000 4800 -2400
rect 5100 -4000 5500 -2400
rect 5800 -4000 6200 -2400
rect 6500 -4000 6900 -2400
rect 7200 -4000 7600 -2400
rect 7900 -4000 8300 -2400
rect 8600 -4000 9000 -2400
rect 9300 -4000 9700 -2400
rect 10000 -4000 10400 -2400
rect 10700 -4000 11100 -2400
<< ndiff >>
rect -2200 1585 -1900 1600
rect -2200 15 -2185 1585
rect -1915 15 -1900 1585
rect -2200 0 -1900 15
rect -1500 1585 -1200 1600
rect -1500 15 -1485 1585
rect -1215 15 -1200 1585
rect -1500 0 -1200 15
rect -800 1585 -500 1600
rect -800 15 -785 1585
rect -515 15 -500 1585
rect -800 0 -500 15
rect -100 1585 200 1600
rect -100 15 -85 1585
rect 185 15 200 1585
rect -100 0 200 15
rect 600 1585 900 1600
rect 600 15 615 1585
rect 885 15 900 1585
rect 600 0 900 15
rect 1300 1585 1600 1600
rect 1300 15 1315 1585
rect 1585 15 1600 1585
rect 1300 0 1600 15
rect 2000 1585 2300 1600
rect 2000 15 2015 1585
rect 2285 15 2300 1585
rect 2000 0 2300 15
rect 2700 1585 3000 1600
rect 2700 15 2715 1585
rect 2985 15 3000 1585
rect 2700 0 3000 15
rect 3400 1585 3700 1600
rect 3400 15 3415 1585
rect 3685 15 3700 1585
rect 3400 0 3700 15
rect 4100 1585 4400 1600
rect 4100 15 4115 1585
rect 4385 15 4400 1585
rect 4100 0 4400 15
rect 4800 1585 5100 1600
rect 4800 15 4815 1585
rect 5085 15 5100 1585
rect 4800 0 5100 15
rect 5500 1585 5800 1600
rect 5500 15 5515 1585
rect 5785 15 5800 1585
rect 5500 0 5800 15
rect 6200 1585 6500 1600
rect 6200 15 6215 1585
rect 6485 15 6500 1585
rect 6200 0 6500 15
rect 6900 1585 7200 1600
rect 6900 15 6915 1585
rect 7185 15 7200 1585
rect 6900 0 7200 15
rect 7600 1585 7900 1600
rect 7600 15 7615 1585
rect 7885 15 7900 1585
rect 7600 0 7900 15
rect 8300 1585 8600 1600
rect 8300 15 8315 1585
rect 8585 15 8600 1585
rect 8300 0 8600 15
rect 9000 1585 9300 1600
rect 9000 15 9015 1585
rect 9285 15 9300 1585
rect 9000 0 9300 15
rect 9700 1585 10000 1600
rect 9700 15 9715 1585
rect 9985 15 10000 1585
rect 9700 0 10000 15
rect 10400 1585 10700 1600
rect 10400 15 10415 1585
rect 10685 15 10700 1585
rect 10400 0 10700 15
rect 11100 1585 11400 1600
rect 11100 15 11115 1585
rect 11385 15 11400 1585
rect 11100 0 11400 15
rect -2200 -415 -1900 -400
rect -2200 -1985 -2185 -415
rect -1915 -1985 -1900 -415
rect -2200 -2000 -1900 -1985
rect -1500 -415 -1200 -400
rect -1500 -1985 -1485 -415
rect -1215 -1985 -1200 -415
rect -1500 -2000 -1200 -1985
rect -800 -415 -500 -400
rect -800 -1985 -785 -415
rect -515 -1985 -500 -415
rect -800 -2000 -500 -1985
rect -100 -415 200 -400
rect -100 -1985 -85 -415
rect 185 -1985 200 -415
rect -100 -2000 200 -1985
rect 600 -415 900 -400
rect 600 -1985 615 -415
rect 885 -1985 900 -415
rect 600 -2000 900 -1985
rect 1300 -415 1600 -400
rect 1300 -1985 1315 -415
rect 1585 -1985 1600 -415
rect 1300 -2000 1600 -1985
rect 2000 -415 2300 -400
rect 2000 -1985 2015 -415
rect 2285 -1985 2300 -415
rect 2000 -2000 2300 -1985
rect 2700 -415 3000 -400
rect 2700 -1985 2715 -415
rect 2985 -1985 3000 -415
rect 2700 -2000 3000 -1985
rect 3400 -415 3700 -400
rect 3400 -1985 3415 -415
rect 3685 -1985 3700 -415
rect 3400 -2000 3700 -1985
rect 4100 -415 4400 -400
rect 4100 -1985 4115 -415
rect 4385 -1985 4400 -415
rect 4100 -2000 4400 -1985
rect 4800 -415 5100 -400
rect 4800 -1985 4815 -415
rect 5085 -1985 5100 -415
rect 4800 -2000 5100 -1985
rect 5500 -415 5800 -400
rect 5500 -1985 5515 -415
rect 5785 -1985 5800 -415
rect 5500 -2000 5800 -1985
rect 6200 -415 6500 -400
rect 6200 -1985 6215 -415
rect 6485 -1985 6500 -415
rect 6200 -2000 6500 -1985
rect 6900 -415 7200 -400
rect 6900 -1985 6915 -415
rect 7185 -1985 7200 -415
rect 6900 -2000 7200 -1985
rect 7600 -415 7900 -400
rect 7600 -1985 7615 -415
rect 7885 -1985 7900 -415
rect 7600 -2000 7900 -1985
rect 8300 -415 8600 -400
rect 8300 -1985 8315 -415
rect 8585 -1985 8600 -415
rect 8300 -2000 8600 -1985
rect 9000 -415 9300 -400
rect 9000 -1985 9015 -415
rect 9285 -1985 9300 -415
rect 9000 -2000 9300 -1985
rect 9700 -415 10000 -400
rect 9700 -1985 9715 -415
rect 9985 -1985 10000 -415
rect 9700 -2000 10000 -1985
rect 10400 -415 10700 -400
rect 10400 -1985 10415 -415
rect 10685 -1985 10700 -415
rect 10400 -2000 10700 -1985
rect 11100 -415 11400 -400
rect 11100 -1985 11115 -415
rect 11385 -1985 11400 -415
rect 11100 -2000 11400 -1985
rect -2200 -2415 -1900 -2400
rect -2200 -3985 -2185 -2415
rect -1915 -3985 -1900 -2415
rect -2200 -4000 -1900 -3985
rect -1500 -2415 -1200 -2400
rect -1500 -3985 -1485 -2415
rect -1215 -3985 -1200 -2415
rect -1500 -4000 -1200 -3985
rect -800 -2415 -500 -2400
rect -800 -3985 -785 -2415
rect -515 -3985 -500 -2415
rect -800 -4000 -500 -3985
rect -100 -2415 200 -2400
rect -100 -3985 -85 -2415
rect 185 -3985 200 -2415
rect -100 -4000 200 -3985
rect 600 -2415 900 -2400
rect 600 -3985 615 -2415
rect 885 -3985 900 -2415
rect 600 -4000 900 -3985
rect 1300 -2415 1600 -2400
rect 1300 -3985 1315 -2415
rect 1585 -3985 1600 -2415
rect 1300 -4000 1600 -3985
rect 2000 -2415 2300 -2400
rect 2000 -3985 2015 -2415
rect 2285 -3985 2300 -2415
rect 2000 -4000 2300 -3985
rect 2700 -2415 3000 -2400
rect 2700 -3985 2715 -2415
rect 2985 -3985 3000 -2415
rect 2700 -4000 3000 -3985
rect 3400 -2415 3700 -2400
rect 3400 -3985 3415 -2415
rect 3685 -3985 3700 -2415
rect 3400 -4000 3700 -3985
rect 4100 -2415 4400 -2400
rect 4100 -3985 4115 -2415
rect 4385 -3985 4400 -2415
rect 4100 -4000 4400 -3985
rect 4800 -2415 5100 -2400
rect 4800 -3985 4815 -2415
rect 5085 -3985 5100 -2415
rect 4800 -4000 5100 -3985
rect 5500 -2415 5800 -2400
rect 5500 -3985 5515 -2415
rect 5785 -3985 5800 -2415
rect 5500 -4000 5800 -3985
rect 6200 -2415 6500 -2400
rect 6200 -3985 6215 -2415
rect 6485 -3985 6500 -2415
rect 6200 -4000 6500 -3985
rect 6900 -2415 7200 -2400
rect 6900 -3985 6915 -2415
rect 7185 -3985 7200 -2415
rect 6900 -4000 7200 -3985
rect 7600 -2415 7900 -2400
rect 7600 -3985 7615 -2415
rect 7885 -3985 7900 -2415
rect 7600 -4000 7900 -3985
rect 8300 -2415 8600 -2400
rect 8300 -3985 8315 -2415
rect 8585 -3985 8600 -2415
rect 8300 -4000 8600 -3985
rect 9000 -2415 9300 -2400
rect 9000 -3985 9015 -2415
rect 9285 -3985 9300 -2415
rect 9000 -4000 9300 -3985
rect 9700 -2415 10000 -2400
rect 9700 -3985 9715 -2415
rect 9985 -3985 10000 -2415
rect 9700 -4000 10000 -3985
rect 10400 -2415 10700 -2400
rect 10400 -3985 10415 -2415
rect 10685 -3985 10700 -2415
rect 10400 -4000 10700 -3985
rect 11100 -2415 11400 -2400
rect 11100 -3985 11115 -2415
rect 11385 -3985 11400 -2415
rect 11100 -4000 11400 -3985
<< ndiffc >>
rect -2185 15 -1915 1585
rect -1485 15 -1215 1585
rect -785 15 -515 1585
rect -85 15 185 1585
rect 615 15 885 1585
rect 1315 15 1585 1585
rect 2015 15 2285 1585
rect 2715 15 2985 1585
rect 3415 15 3685 1585
rect 4115 15 4385 1585
rect 4815 15 5085 1585
rect 5515 15 5785 1585
rect 6215 15 6485 1585
rect 6915 15 7185 1585
rect 7615 15 7885 1585
rect 8315 15 8585 1585
rect 9015 15 9285 1585
rect 9715 15 9985 1585
rect 10415 15 10685 1585
rect 11115 15 11385 1585
rect -2185 -1985 -1915 -415
rect -1485 -1985 -1215 -415
rect -785 -1985 -515 -415
rect -85 -1985 185 -415
rect 615 -1985 885 -415
rect 1315 -1985 1585 -415
rect 2015 -1985 2285 -415
rect 2715 -1985 2985 -415
rect 3415 -1985 3685 -415
rect 4115 -1985 4385 -415
rect 4815 -1985 5085 -415
rect 5515 -1985 5785 -415
rect 6215 -1985 6485 -415
rect 6915 -1985 7185 -415
rect 7615 -1985 7885 -415
rect 8315 -1985 8585 -415
rect 9015 -1985 9285 -415
rect 9715 -1985 9985 -415
rect 10415 -1985 10685 -415
rect 11115 -1985 11385 -415
rect -2185 -3985 -1915 -2415
rect -1485 -3985 -1215 -2415
rect -785 -3985 -515 -2415
rect -85 -3985 185 -2415
rect 615 -3985 885 -2415
rect 1315 -3985 1585 -2415
rect 2015 -3985 2285 -2415
rect 2715 -3985 2985 -2415
rect 3415 -3985 3685 -2415
rect 4115 -3985 4385 -2415
rect 4815 -3985 5085 -2415
rect 5515 -3985 5785 -2415
rect 6215 -3985 6485 -2415
rect 6915 -3985 7185 -2415
rect 7615 -3985 7885 -2415
rect 8315 -3985 8585 -2415
rect 9015 -3985 9285 -2415
rect 9715 -3985 9985 -2415
rect 10415 -3985 10685 -2415
rect 11115 -3985 11385 -2415
<< psubdiff >>
rect 725 1755 775 1770
rect 725 1735 740 1755
rect 760 1735 775 1755
rect 725 1720 775 1735
rect 1425 1725 1475 1740
rect 1425 1705 1440 1725
rect 1460 1705 1475 1725
rect 1425 1690 1475 1705
rect 3525 1730 3575 1745
rect 3525 1710 3540 1730
rect 3560 1710 3575 1730
rect 3525 1695 3575 1710
rect 4225 1725 4275 1740
rect 4225 1705 4240 1725
rect 4260 1705 4275 1725
rect 4225 1690 4275 1705
rect 5625 1730 5675 1745
rect 5625 1710 5640 1730
rect 5660 1710 5675 1730
rect 5625 1695 5675 1710
rect 7025 1725 7075 1740
rect 7025 1705 7040 1725
rect 7060 1705 7075 1725
rect 7025 1690 7075 1705
rect 8425 1725 8475 1740
rect 8425 1705 8440 1725
rect 8460 1705 8475 1725
rect 8425 1690 8475 1705
rect -2500 1585 -2200 1600
rect -2500 15 -2485 1585
rect -2215 15 -2200 1585
rect -2500 0 -2200 15
rect 11400 1585 11700 1600
rect 11400 15 11415 1585
rect 11685 15 11700 1585
rect 11400 0 11700 15
rect 725 -155 775 -140
rect 725 -175 740 -155
rect 760 -175 775 -155
rect 725 -190 775 -175
rect 2825 -235 2875 -220
rect 2825 -255 2840 -235
rect 2860 -255 2875 -235
rect 2825 -270 2875 -255
rect 4925 -235 4975 -220
rect 4925 -255 4940 -235
rect 4960 -255 4975 -235
rect 4925 -270 4975 -255
rect 7725 -205 7775 -190
rect 7725 -225 7740 -205
rect 7760 -225 7775 -205
rect 7725 -240 7775 -225
rect 9125 -235 9175 -220
rect 9125 -255 9140 -235
rect 9160 -255 9175 -235
rect 9125 -270 9175 -255
rect -2500 -415 -2200 -400
rect -2500 -1985 -2485 -415
rect -2215 -1985 -2200 -415
rect -2500 -2000 -2200 -1985
rect 11400 -415 11700 -400
rect 11400 -1985 11415 -415
rect 11685 -1985 11700 -415
rect 11400 -2000 11700 -1985
rect 25 -2335 75 -2320
rect 25 -2355 40 -2335
rect 60 -2355 75 -2335
rect 25 -2370 75 -2355
rect 2825 -2335 2875 -2320
rect 2825 -2355 2840 -2335
rect 2860 -2355 2875 -2335
rect 2825 -2370 2875 -2355
rect 4925 -2330 4975 -2315
rect 4925 -2350 4940 -2330
rect 4960 -2350 4975 -2330
rect 4925 -2365 4975 -2350
rect 7055 -2330 7105 -2315
rect 7055 -2350 7070 -2330
rect 7090 -2350 7105 -2330
rect 7055 -2365 7105 -2350
rect 9125 -2330 9175 -2315
rect 9125 -2350 9140 -2330
rect 9160 -2350 9175 -2330
rect 9125 -2365 9175 -2350
rect -2500 -2415 -2200 -2400
rect -2500 -3985 -2485 -2415
rect -2215 -3985 -2200 -2415
rect -2500 -4000 -2200 -3985
rect 11400 -2415 11700 -2400
rect 11400 -3985 11415 -2415
rect 11685 -3985 11700 -2415
rect 11400 -4000 11700 -3985
rect 725 -4045 775 -4030
rect 725 -4065 740 -4045
rect 760 -4065 775 -4045
rect 2825 -4045 2875 -4030
rect 2825 -4065 2840 -4045
rect 2860 -4065 2875 -4045
rect 4925 -4045 4975 -4030
rect 4925 -4065 4940 -4045
rect 4960 -4065 4975 -4045
rect 7025 -4045 7075 -4030
rect 7025 -4065 7040 -4045
rect 7060 -4065 7075 -4045
rect 9000 -4060 9050 -4055
rect 725 -4080 775 -4065
rect 2825 -4080 2875 -4065
rect 4925 -4080 4975 -4065
rect 7025 -4080 7075 -4065
rect 9000 -4080 9015 -4060
rect 9035 -4080 9050 -4060
rect 9000 -4095 9050 -4080
<< psubdiffcont >>
rect 740 1735 760 1755
rect 1440 1705 1460 1725
rect 3540 1710 3560 1730
rect 4240 1705 4260 1725
rect 5640 1710 5660 1730
rect 7040 1705 7060 1725
rect 8440 1705 8460 1725
rect -2485 15 -2215 1585
rect 11415 15 11685 1585
rect 740 -175 760 -155
rect 2840 -255 2860 -235
rect 4940 -255 4960 -235
rect 7740 -225 7760 -205
rect 9140 -255 9160 -235
rect -2485 -1985 -2215 -415
rect 11415 -1985 11685 -415
rect 40 -2355 60 -2335
rect 2840 -2355 2860 -2335
rect 4940 -2350 4960 -2330
rect 7070 -2350 7090 -2330
rect 9140 -2350 9160 -2330
rect -2485 -3985 -2215 -2415
rect 11415 -3985 11685 -2415
rect 740 -4065 760 -4045
rect 2840 -4065 2860 -4045
rect 4940 -4065 4960 -4045
rect 7040 -4065 7060 -4045
rect 9015 -4080 9035 -4060
<< poly >>
rect 9315 1705 9700 1715
rect 9315 1685 9325 1705
rect 9690 1685 9700 1705
rect 9315 1655 9700 1685
rect -2195 1645 -800 1655
rect -2195 1625 -2185 1645
rect -1915 1625 -1485 1645
rect -1215 1625 -800 1645
rect -2195 1615 -800 1625
rect -1900 1600 -1500 1615
rect -1200 1600 -800 1615
rect -500 1640 9700 1655
rect -500 1600 -100 1640
rect 200 1600 600 1640
rect 900 1600 1300 1615
rect 1600 1600 2000 1640
rect 2300 1600 2700 1615
rect 3000 1600 3400 1640
rect 3700 1600 4100 1615
rect 4400 1600 4800 1640
rect 5100 1600 5500 1615
rect 5800 1600 6200 1640
rect 6500 1600 6900 1615
rect 7200 1600 7600 1640
rect 7900 1600 8300 1615
rect 8600 1600 9000 1640
rect 9300 1600 9700 1640
rect 10000 1645 11395 1655
rect 10000 1625 10415 1645
rect 10685 1625 11115 1645
rect 11385 1625 11395 1645
rect 10000 1615 11395 1625
rect 10000 1600 10400 1615
rect 10700 1600 11100 1615
rect -1900 -15 -1500 0
rect -1200 -15 -800 0
rect -500 -305 -100 0
rect 200 -305 600 0
rect 900 -15 1300 0
rect 1130 -25 1170 -15
rect 1130 -45 1140 -25
rect 1160 -45 1170 -25
rect 1130 -55 1170 -45
rect 1600 -305 2000 0
rect 2300 -15 2700 0
rect 2530 -25 2570 -15
rect 2530 -45 2540 -25
rect 2560 -45 2570 -25
rect 2530 -55 2570 -45
rect 2265 -305 2735 -260
rect 3000 -305 3400 0
rect 3700 -15 4100 0
rect 3830 -25 3870 -15
rect 3830 -45 3840 -25
rect 3860 -45 3870 -25
rect 3830 -55 3870 -45
rect 4400 -305 4800 0
rect 5100 -15 5500 0
rect 5800 -15 6200 0
rect 6500 -15 6900 0
rect 5230 -25 5270 -15
rect 5230 -45 5240 -25
rect 5260 -45 5270 -25
rect 5230 -55 5270 -45
rect 6630 -25 6670 -15
rect 6630 -45 6640 -25
rect 6660 -45 6670 -25
rect 6630 -55 6670 -45
rect 5775 -305 6225 -265
rect 7200 -305 7600 0
rect 7900 -15 8300 0
rect 8030 -25 8070 -15
rect 8030 -45 8040 -25
rect 8060 -45 8070 -25
rect 8030 -55 8070 -45
rect 8600 -305 9000 0
rect 9300 -15 9700 0
rect 10000 -15 10400 0
rect 10700 -15 11100 0
rect -500 -345 2305 -305
rect 2695 -345 5815 -305
rect 6185 -345 9000 -305
rect -2195 -355 -800 -345
rect -2195 -375 -2185 -355
rect -1915 -375 -1485 -355
rect -1215 -375 -800 -355
rect -2195 -385 -800 -375
rect -1900 -400 -1500 -385
rect -1200 -400 -800 -385
rect -500 -400 -100 -345
rect 200 -400 600 -345
rect 900 -400 1300 -345
rect 1600 -400 2000 -345
rect 2530 -355 2570 -345
rect 2530 -375 2540 -355
rect 2560 -375 2570 -355
rect 2530 -385 2570 -375
rect 2300 -400 2700 -385
rect 3000 -400 3400 -345
rect 3700 -400 4100 -345
rect 4400 -400 4800 -345
rect 5100 -400 5500 -345
rect 5930 -355 5970 -345
rect 5930 -375 5940 -355
rect 5960 -375 5970 -355
rect 5930 -385 5970 -375
rect 5800 -400 6200 -385
rect 6500 -400 6900 -345
rect 7200 -400 7600 -345
rect 7900 -400 8300 -345
rect 8600 -400 9000 -345
rect 9705 -355 9995 -345
rect 9705 -370 9715 -355
rect 9300 -375 9715 -370
rect 9985 -370 9995 -355
rect 10405 -355 10695 -345
rect 10405 -370 10415 -355
rect 9985 -375 10415 -370
rect 10685 -370 10695 -355
rect 11105 -355 11395 -345
rect 11105 -370 11115 -355
rect 10685 -375 11115 -370
rect 11385 -375 11395 -355
rect 9300 -385 11395 -375
rect 9300 -400 9700 -385
rect 10000 -400 10400 -385
rect 10700 -400 11100 -385
rect -1900 -2015 -1500 -2000
rect -1200 -2015 -800 -2000
rect -500 -2015 -100 -2000
rect 200 -2015 600 -2000
rect 900 -2015 1300 -2000
rect 1600 -2015 2000 -2000
rect 2300 -2015 2700 -2000
rect 3000 -2015 3400 -2000
rect 3700 -2015 4100 -2000
rect 4400 -2015 4800 -2000
rect 5100 -2015 5500 -2000
rect 5800 -2015 6200 -2000
rect 6500 -2015 6900 -2000
rect 7200 -2015 7600 -2000
rect 7900 -2015 8300 -2000
rect 8600 -2015 9000 -2000
rect 9300 -2015 9700 -2000
rect 10000 -2015 10400 -2000
rect 10700 -2015 11100 -2000
rect 135 -2025 175 -2015
rect 135 -2045 145 -2025
rect 165 -2045 175 -2025
rect 135 -2345 175 -2045
rect 3530 -2025 3570 -2015
rect 3530 -2045 3540 -2025
rect 3560 -2045 3570 -2025
rect 135 -2365 145 -2345
rect 165 -2365 175 -2345
rect 135 -2375 175 -2365
rect 3530 -2355 3570 -2045
rect 6925 -2025 6965 -2015
rect 6925 -2045 6935 -2025
rect 6955 -2045 6965 -2025
rect 6925 -2285 6965 -2045
rect 6925 -2305 6935 -2285
rect 6955 -2305 6965 -2285
rect 6925 -2315 6965 -2305
rect 8325 -2025 8365 -2015
rect 8325 -2045 8335 -2025
rect 8355 -2045 8365 -2025
rect 3530 -2375 3540 -2355
rect 3560 -2375 3570 -2355
rect 8325 -2350 8365 -2045
rect 3530 -2385 3570 -2375
rect 8325 -2370 8335 -2350
rect 8355 -2370 8365 -2350
rect 8325 -2380 8365 -2370
rect -1900 -2400 -1500 -2385
rect -1200 -2400 -800 -2385
rect -500 -2400 -100 -2385
rect 200 -2400 600 -2385
rect 900 -2400 1300 -2385
rect 1600 -2400 2000 -2385
rect 2300 -2400 2700 -2385
rect 3000 -2400 3400 -2385
rect 3700 -2400 4100 -2385
rect 4400 -2400 4800 -2385
rect 5100 -2400 5500 -2385
rect 5800 -2400 6200 -2385
rect 6500 -2400 6900 -2385
rect 7200 -2400 7600 -2385
rect 7900 -2400 8300 -2385
rect 8600 -2400 9000 -2385
rect 9300 -2400 9700 -2385
rect 10000 -2400 10400 -2385
rect 10700 -2400 11100 -2385
rect -1900 -4015 -1500 -4000
rect -1200 -4015 -800 -4000
rect -500 -4015 -100 -4000
rect 200 -4015 600 -4000
rect -2195 -4025 600 -4015
rect -2195 -4045 -2185 -4025
rect -1915 -4045 -1485 -4025
rect -1215 -4045 -785 -4025
rect -515 -4045 -85 -4025
rect 185 -4045 600 -4025
rect -2195 -4055 600 -4045
rect 900 -4035 1300 -4000
rect 900 -4055 910 -4035
rect 1290 -4055 1300 -4035
rect 1600 -4025 2000 -4000
rect 1600 -4045 1610 -4025
rect 1990 -4045 2000 -4025
rect 1600 -4055 2000 -4045
rect 2300 -4035 2700 -4000
rect 2300 -4055 2310 -4035
rect 2690 -4055 2700 -4035
rect 900 -4065 1300 -4055
rect 2300 -4065 2700 -4055
rect 3000 -4035 3400 -4000
rect 3000 -4055 3010 -4035
rect 3390 -4055 3400 -4035
rect 3000 -4065 3400 -4055
rect 3700 -4035 4100 -4000
rect 3700 -4055 3710 -4035
rect 4090 -4055 4100 -4035
rect 3700 -4065 4100 -4055
rect 4400 -4035 4800 -4000
rect 4400 -4055 4410 -4035
rect 4790 -4055 4800 -4035
rect 4400 -4065 4800 -4055
rect 5100 -4035 5500 -4000
rect 5100 -4055 5110 -4035
rect 5485 -4055 5500 -4035
rect 5100 -4065 5500 -4055
rect 5800 -4035 6200 -4000
rect 5800 -4055 5805 -4035
rect 6190 -4055 6200 -4035
rect 5800 -4065 6200 -4055
rect 6500 -4035 6900 -4000
rect 6500 -4055 6510 -4035
rect 6890 -4055 6900 -4035
rect 6500 -4065 6900 -4055
rect 7200 -4035 7600 -4000
rect 7200 -4055 7210 -4035
rect 7590 -4055 7600 -4035
rect 7900 -4015 8300 -4000
rect 8600 -4015 9000 -4000
rect 9300 -4015 9700 -4000
rect 10000 -4015 10400 -4000
rect 10700 -4015 11100 -4000
rect 7900 -4025 11395 -4015
rect 7900 -4045 8315 -4025
rect 8585 -4045 9085 -4025
rect 9285 -4045 9715 -4025
rect 9985 -4045 10415 -4025
rect 10685 -4045 11115 -4025
rect 11385 -4045 11395 -4025
rect 7900 -4055 11395 -4045
rect 7200 -4065 7600 -4055
<< polycont >>
rect 9325 1685 9690 1705
rect -2185 1625 -1915 1645
rect -1485 1625 -1215 1645
rect 10415 1625 10685 1645
rect 11115 1625 11385 1645
rect 1140 -45 1160 -25
rect 2540 -45 2560 -25
rect 3840 -45 3860 -25
rect 5240 -45 5260 -25
rect 6640 -45 6660 -25
rect 8040 -45 8060 -25
rect -2185 -375 -1915 -355
rect -1485 -375 -1215 -355
rect 2540 -375 2560 -355
rect 5940 -375 5960 -355
rect 9715 -375 9985 -355
rect 10415 -375 10685 -355
rect 11115 -375 11385 -355
rect 145 -2045 165 -2025
rect 3540 -2045 3560 -2025
rect 145 -2365 165 -2345
rect 6935 -2045 6955 -2025
rect 6935 -2305 6955 -2285
rect 8335 -2045 8355 -2025
rect 3540 -2375 3560 -2355
rect 8335 -2370 8355 -2350
rect -2185 -4045 -1915 -4025
rect -1485 -4045 -1215 -4025
rect -785 -4045 -515 -4025
rect -85 -4045 185 -4025
rect 910 -4055 1290 -4035
rect 1610 -4045 1990 -4025
rect 2310 -4055 2690 -4035
rect 3010 -4055 3390 -4035
rect 3710 -4055 4090 -4035
rect 4410 -4055 4790 -4035
rect 5110 -4055 5485 -4035
rect 5805 -4055 6190 -4035
rect 6510 -4055 6890 -4035
rect 7210 -4055 7590 -4035
rect 8315 -4045 8585 -4025
rect 9085 -4045 9285 -4025
rect 9715 -4045 9985 -4025
rect 10415 -4045 10685 -4025
rect 11115 -4045 11385 -4025
<< locali >>
rect 730 1755 770 1765
rect 730 1735 740 1755
rect 760 1735 770 1755
rect 9005 1740 11700 1780
rect 730 1725 770 1735
rect 1430 1725 1470 1735
rect 1430 1705 1440 1725
rect 1460 1705 1470 1725
rect 1430 1695 1470 1705
rect 3530 1730 3570 1740
rect 3530 1710 3540 1730
rect 3560 1710 3570 1730
rect 3530 1700 3570 1710
rect 4230 1725 4270 1735
rect 4230 1705 4240 1725
rect 4260 1705 4270 1725
rect 4230 1695 4270 1705
rect 5630 1730 5670 1740
rect 5630 1710 5640 1730
rect 5660 1710 5670 1730
rect 5630 1700 5670 1710
rect 7030 1725 7070 1735
rect 7030 1705 7040 1725
rect 7060 1705 7070 1725
rect 7030 1695 7070 1705
rect 8430 1725 8470 1735
rect 8430 1705 8440 1725
rect 8460 1705 8470 1725
rect 8430 1695 8470 1705
rect -2195 1645 -1905 1655
rect -2195 1625 -2185 1645
rect -1915 1625 -1905 1645
rect -2195 1595 -1905 1625
rect -2495 1585 -1905 1595
rect -2495 15 -2485 1585
rect -2215 15 -2185 1585
rect -1915 15 -1905 1585
rect -2495 5 -1905 15
rect -1495 1645 -1205 1655
rect -1495 1625 -1485 1645
rect -1215 1625 -1205 1645
rect -1495 1585 -1205 1625
rect -1495 15 -1485 1585
rect -1215 15 -1205 1585
rect -1495 5 -1205 15
rect -795 1585 -505 1595
rect -795 15 -785 1585
rect -515 15 -505 1585
rect -795 -20 -505 15
rect -95 1585 195 1595
rect -95 15 -85 1585
rect 185 15 195 1585
rect -95 5 195 15
rect 605 1585 900 1595
rect 605 15 615 1585
rect 885 15 900 1585
rect 605 5 900 15
rect 1305 1585 1595 1595
rect 1305 15 1315 1585
rect 1585 15 1595 1585
rect 605 -20 895 5
rect -795 -60 895 -20
rect 1130 -25 1170 -15
rect 1130 -45 1140 -25
rect 1160 -45 1170 -25
rect 1305 -40 1595 15
rect 2005 1585 2295 1595
rect 2005 15 2015 1585
rect 2285 15 2295 1585
rect 2005 5 2295 15
rect 2705 1585 2995 1595
rect 2705 15 2715 1585
rect 2985 15 2995 1585
rect 2705 5 2995 15
rect 3405 1585 3695 1595
rect 3405 15 3415 1585
rect 3685 15 3695 1585
rect 2530 -25 2570 -15
rect 1130 -55 1170 -45
rect -2195 -355 -1905 -345
rect -2195 -375 -2185 -355
rect -1915 -375 -1905 -355
rect -2195 -405 -1905 -375
rect -2495 -415 -1905 -405
rect -2495 -1985 -2485 -415
rect -2215 -1985 -2185 -415
rect -1915 -1985 -1905 -415
rect -2495 -1995 -1905 -1985
rect -1495 -355 -1205 -345
rect -1495 -375 -1485 -355
rect -1215 -375 -1205 -355
rect -1495 -415 -1205 -375
rect -1495 -1985 -1485 -415
rect -1215 -1985 -1205 -415
rect -1495 -1995 -1205 -1985
rect -795 -415 -505 -405
rect -795 -1985 -785 -415
rect -515 -1985 -505 -415
rect -795 -2080 -505 -1985
rect -95 -415 195 -60
rect 730 -155 770 -145
rect 730 -175 740 -155
rect 760 -175 770 -155
rect 730 -185 770 -175
rect 1420 -255 1460 -40
rect 2530 -45 2540 -25
rect 2560 -45 2570 -25
rect 2530 -55 2570 -45
rect -95 -1985 -85 -415
rect 185 -1985 195 -415
rect -95 -2015 195 -1985
rect 605 -295 1460 -255
rect 2830 -235 2870 -220
rect 2830 -255 2840 -235
rect 2860 -255 2870 -235
rect 2830 -265 2870 -255
rect 605 -405 895 -295
rect 2280 -320 2720 -280
rect 3405 -320 3695 15
rect 4105 1585 4395 1595
rect 4105 15 4115 1585
rect 4385 15 4395 1585
rect 3830 -25 3870 -15
rect 3830 -45 3840 -25
rect 3860 -45 3870 -25
rect 3830 -55 3870 -45
rect 1305 -360 2320 -320
rect 2530 -355 2570 -345
rect 605 -415 900 -405
rect 605 -1985 615 -415
rect 885 -1985 900 -415
rect 605 -1995 900 -1985
rect 1305 -415 1595 -360
rect 2530 -375 2540 -355
rect 2560 -375 2570 -355
rect 2680 -360 3695 -320
rect 2530 -385 2570 -375
rect 1305 -1985 1315 -415
rect 1585 -1985 1595 -415
rect 1305 -1995 1595 -1985
rect 2005 -415 2295 -405
rect 2005 -1985 2015 -415
rect 2285 -1985 2295 -415
rect 135 -2025 175 -2015
rect 135 -2045 145 -2025
rect 165 -2045 175 -2025
rect 135 -2055 175 -2045
rect 605 -2080 895 -1995
rect 2005 -2080 2295 -1985
rect -795 -2120 2295 -2080
rect 2705 -415 2995 -405
rect 2705 -1985 2715 -415
rect 2985 -1985 2995 -415
rect 2705 -2080 2995 -1985
rect 3405 -415 3695 -360
rect 3405 -1985 3415 -415
rect 3685 -1985 3695 -415
rect 3405 -2015 3695 -1985
rect 4105 -320 4395 15
rect 4805 1585 5095 1595
rect 4805 15 4815 1585
rect 5085 15 5095 1585
rect 4805 5 5095 15
rect 5505 1585 5795 1595
rect 5505 15 5515 1585
rect 5785 15 5795 1585
rect 5230 -25 5270 -15
rect 5230 -45 5240 -25
rect 5260 -45 5270 -25
rect 5230 -55 5270 -45
rect 4930 -235 4970 -225
rect 4930 -255 4940 -235
rect 4960 -255 4970 -235
rect 4930 -265 4970 -255
rect 5505 -260 5795 15
rect 6205 1585 6495 1595
rect 6205 15 6215 1585
rect 6485 15 6495 1585
rect 6205 5 6495 15
rect 6905 1585 7195 1595
rect 6905 15 6915 1585
rect 7185 15 7195 1585
rect 6630 -25 6670 -15
rect 6630 -45 6640 -25
rect 6660 -45 6670 -25
rect 6630 -55 6670 -45
rect 6905 -260 7195 15
rect 7605 1585 7895 1595
rect 7605 15 7615 1585
rect 7885 15 7895 1585
rect 7605 5 7895 15
rect 8305 1585 8595 1595
rect 8305 15 8315 1585
rect 8585 15 8595 1585
rect 8030 -25 8070 -15
rect 8030 -45 8040 -25
rect 8060 -45 8070 -25
rect 8030 -55 8070 -45
rect 8305 -20 8595 15
rect 9005 1585 9295 1740
rect 9315 1705 11700 1715
rect 9315 1685 9325 1705
rect 9690 1685 11700 1705
rect 9315 1675 11700 1685
rect 10405 1645 10695 1655
rect 10405 1625 10415 1645
rect 10685 1625 10695 1645
rect 9005 15 9015 1585
rect 9285 15 9295 1585
rect 9005 5 9295 15
rect 9705 1585 9995 1595
rect 9705 15 9715 1585
rect 9985 15 9995 1585
rect 9705 -20 9995 15
rect 10405 1585 10695 1625
rect 10405 15 10415 1585
rect 10685 15 10695 1585
rect 10405 5 10695 15
rect 11105 1645 11395 1655
rect 11105 1625 11115 1645
rect 11385 1625 11395 1645
rect 11105 1595 11395 1625
rect 11105 1585 11695 1595
rect 11105 15 11115 1585
rect 11385 15 11415 1585
rect 11685 15 11695 1585
rect 11105 5 11695 15
rect 8305 -60 9995 -20
rect 7730 -205 7770 -195
rect 7730 -225 7740 -205
rect 7760 -225 7770 -205
rect 7730 -235 7770 -225
rect 5505 -300 6220 -260
rect 6905 -300 7895 -260
rect 6180 -320 6220 -300
rect 4105 -360 5795 -320
rect 4105 -415 4395 -360
rect 4105 -1985 4115 -415
rect 4385 -1985 4395 -415
rect 3530 -2025 3570 -2015
rect 3530 -2045 3540 -2025
rect 3560 -2045 3570 -2025
rect 3530 -2055 3570 -2045
rect 4105 -2080 4395 -1985
rect 4805 -415 5095 -405
rect 4805 -1985 4815 -415
rect 5085 -1985 5095 -415
rect 4805 -2015 5095 -1985
rect 5505 -415 5795 -360
rect 5930 -355 5970 -345
rect 5930 -375 5940 -355
rect 5960 -375 5970 -355
rect 6180 -360 7195 -320
rect 5930 -385 5970 -375
rect 5505 -1985 5515 -415
rect 5785 -1985 5795 -415
rect 5505 -1995 5795 -1985
rect 6205 -415 6495 -405
rect 6205 -1985 6215 -415
rect 6485 -1985 6495 -415
rect 2705 -2120 4395 -2080
rect 30 -2335 70 -2325
rect 30 -2355 40 -2335
rect 60 -2355 70 -2335
rect 30 -2405 70 -2355
rect 135 -2345 1595 -2335
rect 135 -2365 145 -2345
rect 165 -2365 1595 -2345
rect 135 -2375 1595 -2365
rect -2495 -2415 -1905 -2405
rect -2495 -3985 -2485 -2415
rect -2215 -3985 -2185 -2415
rect -1915 -3985 -1905 -2415
rect -2495 -3995 -1905 -3985
rect -2195 -4025 -1905 -3995
rect -2195 -4045 -2185 -4025
rect -1915 -4045 -1905 -4025
rect -2195 -4055 -1905 -4045
rect -1495 -2415 -1205 -2405
rect -1495 -3985 -1485 -2415
rect -1215 -3985 -1205 -2415
rect -1495 -4025 -1205 -3985
rect -1495 -4045 -1485 -4025
rect -1215 -4045 -1205 -4025
rect -1495 -4055 -1205 -4045
rect -795 -2415 -505 -2405
rect -795 -3985 -785 -2415
rect -515 -3985 -505 -2415
rect -795 -4025 -505 -3985
rect -795 -4045 -785 -4025
rect -515 -4045 -505 -4025
rect -795 -4055 -505 -4045
rect -95 -2415 195 -2405
rect -95 -3985 -85 -2415
rect 185 -3985 195 -2415
rect -95 -4025 195 -3985
rect 605 -2415 900 -2405
rect 605 -3985 615 -2415
rect 885 -3985 900 -2415
rect 605 -3995 900 -3985
rect 1305 -2415 1595 -2375
rect 1305 -3985 1315 -2415
rect 1585 -3985 1595 -2415
rect 1305 -3995 1595 -3985
rect 2005 -2415 2295 -2120
rect 2830 -2335 2870 -2325
rect 2830 -2355 2840 -2335
rect 2860 -2355 2870 -2335
rect 2830 -2405 2870 -2355
rect 3530 -2355 3570 -2345
rect 3530 -2375 3540 -2355
rect 3560 -2375 3570 -2355
rect 3530 -2385 3570 -2375
rect 2005 -3985 2015 -2415
rect 2285 -3985 2295 -2415
rect 2005 -3995 2295 -3985
rect 2705 -2415 2995 -2405
rect 2705 -3985 2715 -2415
rect 2985 -3985 2995 -2415
rect 2705 -3995 2995 -3985
rect 3405 -2415 3695 -2385
rect 3405 -3985 3415 -2415
rect 3685 -3985 3695 -2415
rect 3405 -3995 3695 -3985
rect 4105 -2415 4395 -2120
rect 5055 -2275 5095 -2015
rect 6205 -2080 6495 -1985
rect 6905 -415 7195 -360
rect 6905 -1985 6915 -415
rect 7185 -1985 7195 -415
rect 6905 -2015 7195 -1985
rect 7605 -415 7895 -300
rect 7605 -1985 7615 -415
rect 7885 -1985 7895 -415
rect 6925 -2025 6965 -2015
rect 6925 -2045 6935 -2025
rect 6955 -2045 6965 -2025
rect 6925 -2055 6965 -2045
rect 7605 -2080 7895 -1985
rect 8305 -415 8595 -60
rect 9130 -235 9170 -225
rect 9130 -255 9140 -235
rect 9160 -255 9170 -235
rect 9130 -265 9170 -255
rect 9705 -355 9995 -345
rect 9705 -375 9715 -355
rect 9985 -375 9995 -355
rect 8305 -1985 8315 -415
rect 8585 -1985 8595 -415
rect 8305 -2015 8595 -1985
rect 9005 -415 9295 -405
rect 9005 -1985 9015 -415
rect 9285 -1985 9295 -415
rect 8325 -2025 8365 -2015
rect 8325 -2045 8335 -2025
rect 8355 -2045 8365 -2025
rect 8325 -2055 8365 -2045
rect 9005 -2080 9295 -1985
rect 9705 -415 9995 -375
rect 9705 -1985 9715 -415
rect 9985 -1985 9995 -415
rect 9705 -1995 9995 -1985
rect 10405 -355 10695 -345
rect 10405 -375 10415 -355
rect 10685 -375 10695 -355
rect 10405 -415 10695 -375
rect 10405 -1985 10415 -415
rect 10685 -1985 10695 -415
rect 10405 -1995 10695 -1985
rect 11105 -355 11395 -345
rect 11105 -375 11115 -355
rect 11385 -375 11395 -355
rect 11105 -405 11395 -375
rect 11105 -415 11695 -405
rect 11105 -1985 11115 -415
rect 11385 -1985 11415 -415
rect 11685 -1985 11695 -415
rect 11105 -1995 11695 -1985
rect 6205 -2120 9295 -2080
rect 5055 -2285 6965 -2275
rect 5055 -2305 6935 -2285
rect 6955 -2305 6965 -2285
rect 5055 -2315 6965 -2305
rect 4930 -2330 4970 -2320
rect 4930 -2350 4940 -2330
rect 4960 -2350 4970 -2330
rect 4930 -2405 4970 -2350
rect 4105 -3985 4115 -2415
rect 4385 -3985 4395 -2415
rect 4105 -3995 4395 -3985
rect 4805 -2415 5095 -2405
rect 4805 -3985 4815 -2415
rect 5085 -3985 5095 -2415
rect 4805 -3995 5095 -3985
rect 5505 -2415 5795 -2315
rect 6985 -2340 7025 -2120
rect 5505 -3985 5515 -2415
rect 5785 -3985 5795 -2415
rect 5505 -3995 5795 -3985
rect 6205 -2380 7025 -2340
rect 7060 -2330 7100 -2320
rect 7060 -2350 7070 -2330
rect 7090 -2350 7100 -2330
rect 9130 -2330 9170 -2320
rect 6205 -2415 6495 -2380
rect 7060 -2405 7100 -2350
rect 8325 -2350 8365 -2340
rect 8325 -2360 8335 -2350
rect 7605 -2370 8335 -2360
rect 8355 -2370 8365 -2350
rect 7605 -2380 8365 -2370
rect 9130 -2350 9140 -2330
rect 9160 -2350 9170 -2330
rect 6205 -3985 6215 -2415
rect 6485 -3985 6495 -2415
rect 6205 -3995 6495 -3985
rect 6905 -2415 7195 -2405
rect 6905 -3985 6915 -2415
rect 7185 -3985 7195 -2415
rect 6905 -3995 7195 -3985
rect 7605 -2415 7895 -2380
rect 9130 -2405 9170 -2350
rect 7605 -3985 7615 -2415
rect 7885 -3985 7895 -2415
rect 7605 -3995 7895 -3985
rect 8305 -2415 8595 -2405
rect 8305 -3985 8315 -2415
rect 8585 -3985 8595 -2415
rect -95 -4045 -85 -4025
rect 185 -4045 195 -4025
rect -95 -4055 195 -4045
rect 730 -4045 770 -3995
rect 1600 -4025 2000 -4015
rect 730 -4065 740 -4045
rect 760 -4065 770 -4045
rect 900 -4035 1300 -4025
rect 900 -4055 910 -4035
rect 1290 -4055 1300 -4035
rect 1600 -4045 1610 -4025
rect 1990 -4045 2000 -4025
rect 1600 -4055 2000 -4045
rect 2300 -4035 2700 -4025
rect 2300 -4055 2310 -4035
rect 2690 -4055 2700 -4035
rect 900 -4065 1300 -4055
rect 2300 -4065 2700 -4055
rect 2830 -4045 2870 -3995
rect 2830 -4065 2840 -4045
rect 2860 -4065 2870 -4045
rect 3000 -4035 3400 -4025
rect 3000 -4055 3010 -4035
rect 3390 -4055 3400 -4035
rect 3000 -4065 3400 -4055
rect 3700 -4035 4100 -4025
rect 3700 -4055 3710 -4035
rect 4090 -4055 4100 -4035
rect 3700 -4065 4100 -4055
rect 4400 -4035 4800 -4025
rect 4400 -4055 4410 -4035
rect 4790 -4055 4800 -4035
rect 4400 -4065 4800 -4055
rect 4930 -4045 4970 -3995
rect 4930 -4065 4940 -4045
rect 4960 -4065 4970 -4045
rect 5100 -4035 5495 -4025
rect 5100 -4055 5110 -4035
rect 5485 -4055 5495 -4035
rect 5100 -4065 5495 -4055
rect 5800 -4035 6200 -4025
rect 5800 -4055 5805 -4035
rect 6190 -4055 6200 -4035
rect 5800 -4065 6200 -4055
rect 6500 -4035 6900 -4025
rect 6500 -4055 6510 -4035
rect 6890 -4055 6900 -4035
rect 6500 -4065 6900 -4055
rect 7030 -4045 7070 -3995
rect 8305 -4025 8595 -3985
rect 7030 -4065 7040 -4045
rect 7060 -4065 7070 -4045
rect 7200 -4035 7600 -4025
rect 7200 -4055 7210 -4035
rect 7590 -4055 7600 -4035
rect 8305 -4045 8315 -4025
rect 8585 -4045 8595 -4025
rect 8305 -4055 8595 -4045
rect 9005 -2415 9295 -2405
rect 9005 -3985 9015 -2415
rect 9285 -3985 9295 -2415
rect 9005 -4015 9295 -3985
rect 7200 -4065 7600 -4055
rect 9005 -4060 9045 -4015
rect 9075 -4025 9295 -4015
rect 9075 -4045 9085 -4025
rect 9285 -4045 9295 -4025
rect 9075 -4055 9295 -4045
rect 9705 -2415 9995 -2405
rect 9705 -3985 9715 -2415
rect 9985 -3985 9995 -2415
rect 9705 -4025 9995 -3985
rect 9705 -4045 9715 -4025
rect 9985 -4045 9995 -4025
rect 9705 -4055 9995 -4045
rect 10405 -2415 10695 -2405
rect 10405 -3985 10415 -2415
rect 10685 -3985 10695 -2415
rect 10405 -4025 10695 -3985
rect 10405 -4045 10415 -4025
rect 10685 -4045 10695 -4025
rect 10405 -4055 10695 -4045
rect 11105 -2415 11695 -2405
rect 11105 -3985 11115 -2415
rect 11385 -3985 11415 -2415
rect 11685 -3985 11695 -2415
rect 11105 -3995 11695 -3985
rect 11105 -4025 11395 -3995
rect 11105 -4045 11115 -4025
rect 11385 -4045 11395 -4025
rect 11105 -4055 11395 -4045
rect 730 -4075 770 -4065
rect 2830 -4075 2870 -4065
rect 4930 -4075 4970 -4065
rect 7030 -4075 7070 -4065
rect 9005 -4080 9015 -4060
rect 9035 -4080 9045 -4060
rect 9005 -4090 9045 -4080
<< viali >>
rect 740 1735 760 1755
rect 1440 1705 1460 1725
rect 3540 1710 3560 1730
rect 4240 1705 4260 1725
rect 5640 1710 5660 1730
rect 7040 1705 7060 1725
rect 8440 1705 8460 1725
rect -2485 15 -2215 1585
rect -2185 15 -1915 1585
rect -1485 15 -1215 1585
rect -85 15 185 1585
rect 1140 -45 1160 -25
rect 2015 15 2285 1585
rect 2715 15 2985 1585
rect -2485 -1985 -2215 -415
rect -2185 -1985 -1915 -415
rect -1485 -1985 -1215 -415
rect 740 -175 760 -155
rect 2540 -45 2560 -25
rect 2840 -255 2860 -235
rect 3840 -45 3860 -25
rect 2540 -375 2560 -355
rect 4815 15 5085 1585
rect 5240 -45 5260 -25
rect 4940 -255 4960 -235
rect 6215 15 6485 1585
rect 6640 -45 6660 -25
rect 7615 15 7885 1585
rect 8040 -45 8060 -25
rect 10415 15 10685 1585
rect 11115 15 11385 1585
rect 11415 15 11685 1585
rect 7740 -225 7760 -205
rect 5940 -375 5960 -355
rect -2485 -3985 -2215 -2415
rect -2185 -3985 -1915 -2415
rect -1485 -3985 -1215 -2415
rect -785 -3985 -515 -2415
rect -85 -3985 185 -2415
rect 615 -3985 885 -2415
rect 2715 -3985 2985 -2415
rect 9140 -255 9160 -235
rect 9715 -1985 9985 -415
rect 10415 -1985 10685 -415
rect 11115 -1985 11385 -415
rect 11415 -1985 11685 -415
rect 4815 -3985 5085 -2415
rect 6915 -3985 7185 -2415
rect 8315 -3985 8585 -2415
rect 910 -4055 1290 -4035
rect 1610 -4045 1990 -4025
rect 2310 -4055 2690 -4035
rect 3010 -4055 3390 -4035
rect 3710 -4055 4090 -4035
rect 4410 -4055 4790 -4035
rect 5110 -4055 5485 -4035
rect 5805 -4055 6190 -4035
rect 6510 -4055 6890 -4035
rect 7210 -4055 7590 -4035
rect 9015 -3985 9285 -2415
rect 9715 -3985 9985 -2415
rect 10415 -3985 10685 -2415
rect 11115 -3985 11385 -2415
rect 11415 -3985 11685 -2415
<< metal1 >>
rect -2500 1815 11700 3405
rect -2500 1585 -1205 1595
rect -2500 15 -2485 1585
rect -2215 15 -2185 1585
rect -1915 15 -1485 1585
rect -1215 15 -1205 1585
rect -2500 -400 -1205 15
rect -95 1585 195 1815
rect 725 1755 775 1770
rect 725 1735 740 1755
rect 760 1735 775 1755
rect 725 1690 775 1735
rect 1425 1725 1475 1740
rect 1425 1705 1440 1725
rect 1460 1705 1475 1725
rect 1425 1690 1475 1705
rect -95 15 -85 1585
rect 185 15 195 1585
rect -95 5 195 15
rect 605 -155 895 1690
rect 605 -175 740 -155
rect 760 -175 895 -155
rect 605 -400 895 -175
rect 1130 -25 1170 -15
rect 1130 -45 1140 -25
rect 1160 -45 1170 -25
rect 1130 -400 1170 -45
rect 1305 -400 1595 1690
rect 2005 1585 2295 1815
rect 2005 15 2015 1585
rect 2285 15 2295 1585
rect 2005 5 2295 15
rect 2705 1585 2995 1815
rect 3525 1730 3575 1745
rect 3405 1710 3540 1730
rect 3560 1710 3695 1730
rect 3405 1600 3695 1710
rect 4225 1725 4275 1740
rect 4225 1705 4240 1725
rect 4260 1705 4275 1725
rect 4225 1690 4275 1705
rect 4105 1600 4395 1690
rect 2705 15 2715 1585
rect 2985 15 2995 1585
rect 4805 1585 5095 1815
rect 5625 1730 5675 1745
rect 5625 1710 5640 1730
rect 5660 1710 5675 1730
rect 5625 1690 5675 1710
rect 2705 5 2995 15
rect 2530 -25 2570 -15
rect 2530 -45 2540 -25
rect 2560 -45 2570 -25
rect 2530 -355 2570 -45
rect 2530 -375 2540 -355
rect 2560 -375 2570 -355
rect 2530 -400 2570 -375
rect 2705 -235 2995 -210
rect 2705 -255 2840 -235
rect 2860 -255 2995 -235
rect 2705 -400 2995 -255
rect 3405 -400 3695 1565
rect 3830 -25 3870 -15
rect 3830 -45 3840 -25
rect 3860 -45 3870 -25
rect 3830 -400 3870 -45
rect 4105 -320 4395 1570
rect 4805 15 4815 1585
rect 5085 15 5095 1585
rect 4805 5 5095 15
rect 5230 -25 5270 -15
rect 5230 -45 5240 -25
rect 5260 -45 5270 -25
rect 4805 -235 5095 -210
rect 4805 -255 4940 -235
rect 4960 -255 5095 -235
rect 4805 -320 5095 -255
rect 5230 -320 5270 -45
rect 5505 -320 5795 1690
rect 6205 1585 6495 1815
rect 7025 1725 7075 1740
rect 7025 1705 7040 1725
rect 7060 1705 7075 1725
rect 7025 1690 7075 1705
rect 6205 15 6215 1585
rect 6485 15 6495 1585
rect 6205 5 6495 15
rect 4105 -340 5795 -320
rect 4105 -400 4395 -340
rect 4805 -400 5095 -340
rect 5230 -400 5270 -340
rect 5505 -400 5795 -340
rect 6630 -25 6670 -15
rect 6630 -45 6640 -25
rect 6660 -45 6670 -25
rect 5930 -355 5970 -345
rect 5930 -375 5940 -355
rect 5960 -375 5970 -355
rect 5930 -400 5970 -375
rect 6630 -400 6670 -45
rect 6905 -320 7195 1690
rect 7605 1585 7895 1815
rect 8425 1725 8475 1740
rect 8425 1705 8440 1725
rect 8460 1705 8475 1725
rect 8425 1690 8475 1705
rect 7605 15 7615 1585
rect 7885 15 7895 1585
rect 7605 5 7895 15
rect 8030 -25 8070 -15
rect 8030 -45 8040 -25
rect 8060 -45 8070 -25
rect 6885 -340 7195 -320
rect 6905 -400 7195 -340
rect 7605 -205 7895 -170
rect 7605 -225 7740 -205
rect 7760 -225 7895 -205
rect 7605 -400 7895 -225
rect 8030 -400 8070 -45
rect 8305 -400 8595 1690
rect 10405 1585 11695 1595
rect 10405 15 10415 1585
rect 10685 15 11115 1585
rect 11385 15 11415 1585
rect 11685 15 11695 1585
rect 9005 -235 9295 -175
rect 9005 -255 9140 -235
rect 9160 -255 9295 -235
rect 9005 -400 9295 -255
rect 10405 -400 11695 15
rect -2500 -415 11700 -400
rect -2500 -1985 -2485 -415
rect -2215 -1985 -2185 -415
rect -1915 -1985 -1485 -415
rect -1215 -1985 9715 -415
rect 9985 -1985 10415 -415
rect 10685 -1985 11115 -415
rect 11385 -1985 11415 -415
rect 11685 -1985 11700 -415
rect -2500 -2415 11700 -1985
rect -2500 -3985 -2485 -2415
rect -2215 -3985 -2185 -2415
rect -1915 -3985 -1485 -2415
rect -1215 -3985 -785 -2415
rect -515 -3985 -85 -2415
rect 185 -3985 615 -2415
rect 885 -3985 2715 -2415
rect 2985 -3985 4815 -2415
rect 5085 -3985 6915 -2415
rect 7185 -3985 8315 -2415
rect 8585 -3985 9015 -2415
rect 9285 -3985 9715 -2415
rect 9985 -3985 10415 -2415
rect 10685 -3985 11115 -2415
rect 11385 -3985 11415 -2415
rect 11685 -3985 11700 -2415
rect -2500 -3995 11700 -3985
rect 1600 -4025 2000 -3995
rect 900 -4035 1300 -4025
rect 900 -4055 910 -4035
rect 1290 -4055 1300 -4035
rect 1600 -4045 1610 -4025
rect 1990 -4045 2000 -4025
rect 1600 -4055 2000 -4045
rect 2300 -4035 2700 -4025
rect 2300 -4055 2310 -4035
rect 2690 -4055 2700 -4035
rect 900 -4065 1300 -4055
rect 2300 -4065 2700 -4055
rect 3000 -4035 3400 -4025
rect 3000 -4055 3010 -4035
rect 3390 -4055 3400 -4035
rect 3000 -4065 3400 -4055
rect 3700 -4035 4100 -3995
rect 3700 -4055 3710 -4035
rect 4090 -4055 4100 -4035
rect 3700 -4065 4100 -4055
rect 4400 -4035 4800 -4025
rect 4400 -4055 4410 -4035
rect 4790 -4055 4800 -4035
rect 4400 -4065 4800 -4055
rect 5100 -4035 5500 -4025
rect 5100 -4055 5110 -4035
rect 5485 -4055 5500 -4035
rect 5100 -4065 5500 -4055
rect 5800 -4035 6200 -3995
rect 5800 -4055 5805 -4035
rect 6190 -4055 6200 -4035
rect 5800 -4065 6200 -4055
rect 6500 -4035 6900 -4025
rect 6500 -4055 6510 -4035
rect 6890 -4055 6900 -4035
rect 6500 -4065 6900 -4055
rect 7200 -4035 7600 -4025
rect 7200 -4055 7210 -4035
rect 7590 -4055 7600 -4035
rect 7200 -4065 7600 -4055
<< labels >>
rlabel locali 11700 1695 11700 1695 3 Vg
rlabel poly 7350 -4065 7350 -4065 5 b6
rlabel poly 6650 -4065 6650 -4065 5 b5
rlabel poly 5245 -4065 5245 -4065 5 b4
rlabel poly 4550 -4065 4550 -4065 5 b3
rlabel poly 3150 -4065 3150 -4065 5 b2
rlabel poly 2550 -4065 2550 -4065 5 b1
rlabel poly 1155 -4065 1155 -4065 5 b0
rlabel metal1 -2500 -2215 -2500 -2215 7 GND
rlabel metal1 -2500 2575 -2500 2575 7 VDD
<< end >>
