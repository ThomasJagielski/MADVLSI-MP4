magic
tech sky130A
timestamp 1617442879
<< nmos >>
rect 0 0 300 1600
rect 600 0 900 1600
rect 1200 0 1500 1600
rect 1800 0 2100 1600
rect 2400 0 2700 1600
rect 3000 0 3300 1600
rect 3600 0 3900 1600
rect 4200 0 4500 1600
rect 4800 0 5100 1600
rect 5400 0 5700 1600
rect 6000 0 6300 1600
rect 6600 0 6900 1600
rect 7200 0 7500 1600
rect 7800 0 8100 1600
rect 8400 0 8700 1600
rect 9000 0 9300 1600
rect 9600 0 9900 1600
rect 10200 0 10500 1600
rect 10800 0 11100 1600
rect 0 -2000 300 -400
rect 600 -2000 900 -400
rect 1200 -2000 1500 -400
rect 1800 -2000 2100 -400
rect 2400 -2000 2700 -400
rect 3000 -2000 3300 -400
rect 3600 -2000 3900 -400
rect 4200 -2000 4500 -400
rect 4800 -2000 5100 -400
rect 5400 -2000 5700 -400
rect 6000 -2000 6300 -400
rect 6600 -2000 6900 -400
rect 7200 -2000 7500 -400
rect 7800 -2000 8100 -400
rect 8400 -2000 8700 -400
rect 9000 -2000 9300 -400
rect 9600 -2000 9900 -400
rect 10200 -2000 10500 -400
rect 10800 -2000 11100 -400
rect 0 -4000 300 -2400
rect 600 -4000 900 -2400
rect 1200 -4000 1500 -2400
rect 1800 -4000 2100 -2400
rect 2400 -4000 2700 -2400
rect 3000 -4000 3300 -2400
rect 3600 -4000 3900 -2400
rect 4200 -4000 4500 -2400
rect 4800 -4000 5100 -2400
rect 5400 -4000 5700 -2400
rect 6000 -4000 6300 -2400
rect 6600 -4000 6900 -2400
rect 7200 -4000 7500 -2400
rect 7800 -4000 8100 -2400
rect 8400 -4000 8700 -2400
rect 9000 -4000 9300 -2400
rect 9600 -4000 9900 -2400
rect 10200 -4000 10500 -2400
rect 10800 -4000 11100 -2400
<< ndiff >>
rect -300 1585 0 1600
rect -300 15 -285 1585
rect -15 15 0 1585
rect -300 0 0 15
rect 300 1585 600 1600
rect 300 15 315 1585
rect 585 15 600 1585
rect 300 0 600 15
rect 900 1585 1200 1600
rect 900 15 915 1585
rect 1185 15 1200 1585
rect 900 0 1200 15
rect 1500 1585 1800 1600
rect 1500 15 1515 1585
rect 1785 15 1800 1585
rect 1500 0 1800 15
rect 2100 1585 2400 1600
rect 2100 15 2115 1585
rect 2385 15 2400 1585
rect 2100 0 2400 15
rect 2700 1585 3000 1600
rect 2700 15 2715 1585
rect 2985 15 3000 1585
rect 2700 0 3000 15
rect 3300 1585 3600 1600
rect 3300 15 3315 1585
rect 3585 15 3600 1585
rect 3300 0 3600 15
rect 3900 1585 4200 1600
rect 3900 15 3915 1585
rect 4185 15 4200 1585
rect 3900 0 4200 15
rect 4500 1585 4800 1600
rect 4500 15 4515 1585
rect 4785 15 4800 1585
rect 4500 0 4800 15
rect 5100 1585 5400 1600
rect 5100 15 5115 1585
rect 5385 15 5400 1585
rect 5100 0 5400 15
rect 5700 1585 6000 1600
rect 5700 15 5715 1585
rect 5985 15 6000 1585
rect 5700 0 6000 15
rect 6300 1585 6600 1600
rect 6300 15 6315 1585
rect 6585 15 6600 1585
rect 6300 0 6600 15
rect 6900 1585 7200 1600
rect 6900 15 6915 1585
rect 7185 15 7200 1585
rect 6900 0 7200 15
rect 7500 1585 7800 1600
rect 7500 15 7515 1585
rect 7785 15 7800 1585
rect 7500 0 7800 15
rect 8100 1585 8400 1600
rect 8100 15 8115 1585
rect 8385 15 8400 1585
rect 8100 0 8400 15
rect 8700 1585 9000 1600
rect 8700 15 8715 1585
rect 8985 15 9000 1585
rect 8700 0 9000 15
rect 9300 1585 9600 1600
rect 9300 15 9315 1585
rect 9585 15 9600 1585
rect 9300 0 9600 15
rect 9900 1585 10200 1600
rect 9900 15 9915 1585
rect 10185 15 10200 1585
rect 9900 0 10200 15
rect 10500 1585 10800 1600
rect 10500 15 10515 1585
rect 10785 15 10800 1585
rect 10500 0 10800 15
rect 11100 1585 11400 1600
rect 11100 15 11115 1585
rect 11385 15 11400 1585
rect 11100 0 11400 15
rect -300 -415 0 -400
rect -300 -1985 -285 -415
rect -15 -1985 0 -415
rect -300 -2000 0 -1985
rect 300 -415 600 -400
rect 300 -1985 315 -415
rect 585 -1985 600 -415
rect 300 -2000 600 -1985
rect 900 -415 1200 -400
rect 900 -1985 915 -415
rect 1185 -1985 1200 -415
rect 900 -2000 1200 -1985
rect 1500 -415 1800 -400
rect 1500 -1985 1515 -415
rect 1785 -1985 1800 -415
rect 1500 -2000 1800 -1985
rect 2100 -415 2400 -400
rect 2100 -1985 2115 -415
rect 2385 -1985 2400 -415
rect 2100 -2000 2400 -1985
rect 2700 -415 3000 -400
rect 2700 -1985 2715 -415
rect 2985 -1985 3000 -415
rect 2700 -2000 3000 -1985
rect 3300 -415 3600 -400
rect 3300 -1985 3315 -415
rect 3585 -1985 3600 -415
rect 3300 -2000 3600 -1985
rect 3900 -415 4200 -400
rect 3900 -1985 3915 -415
rect 4185 -1985 4200 -415
rect 3900 -2000 4200 -1985
rect 4500 -415 4800 -400
rect 4500 -1985 4515 -415
rect 4785 -1985 4800 -415
rect 4500 -2000 4800 -1985
rect 5100 -415 5400 -400
rect 5100 -1985 5115 -415
rect 5385 -1985 5400 -415
rect 5100 -2000 5400 -1985
rect 5700 -415 6000 -400
rect 5700 -1985 5715 -415
rect 5985 -1985 6000 -415
rect 5700 -2000 6000 -1985
rect 6300 -415 6600 -400
rect 6300 -1985 6315 -415
rect 6585 -1985 6600 -415
rect 6300 -2000 6600 -1985
rect 6900 -415 7200 -400
rect 6900 -1985 6915 -415
rect 7185 -1985 7200 -415
rect 6900 -2000 7200 -1985
rect 7500 -415 7800 -400
rect 7500 -1985 7515 -415
rect 7785 -1985 7800 -415
rect 7500 -2000 7800 -1985
rect 8100 -415 8400 -400
rect 8100 -1985 8115 -415
rect 8385 -1985 8400 -415
rect 8100 -2000 8400 -1985
rect 8700 -415 9000 -400
rect 8700 -1985 8715 -415
rect 8985 -1985 9000 -415
rect 8700 -2000 9000 -1985
rect 9300 -415 9600 -400
rect 9300 -1985 9315 -415
rect 9585 -1985 9600 -415
rect 9300 -2000 9600 -1985
rect 9900 -415 10200 -400
rect 9900 -1985 9915 -415
rect 10185 -1985 10200 -415
rect 9900 -2000 10200 -1985
rect 10500 -415 10800 -400
rect 10500 -1985 10515 -415
rect 10785 -1985 10800 -415
rect 10500 -2000 10800 -1985
rect 11100 -415 11400 -400
rect 11100 -1985 11115 -415
rect 11385 -1985 11400 -415
rect 11100 -2000 11400 -1985
rect -300 -2415 0 -2400
rect -300 -3985 -285 -2415
rect -15 -3985 0 -2415
rect -300 -4000 0 -3985
rect 300 -2415 600 -2400
rect 300 -3985 315 -2415
rect 585 -3985 600 -2415
rect 300 -4000 600 -3985
rect 900 -2415 1200 -2400
rect 900 -3985 915 -2415
rect 1185 -3985 1200 -2415
rect 900 -4000 1200 -3985
rect 1500 -2415 1800 -2400
rect 1500 -3985 1515 -2415
rect 1785 -3985 1800 -2415
rect 1500 -4000 1800 -3985
rect 2100 -2415 2400 -2400
rect 2100 -3985 2115 -2415
rect 2385 -3985 2400 -2415
rect 2100 -4000 2400 -3985
rect 2700 -2415 3000 -2400
rect 2700 -3985 2715 -2415
rect 2985 -3985 3000 -2415
rect 2700 -4000 3000 -3985
rect 3300 -2415 3600 -2400
rect 3300 -3985 3315 -2415
rect 3585 -3985 3600 -2415
rect 3300 -4000 3600 -3985
rect 3900 -2415 4200 -2400
rect 3900 -3985 3915 -2415
rect 4185 -3985 4200 -2415
rect 3900 -4000 4200 -3985
rect 4500 -2415 4800 -2400
rect 4500 -3985 4515 -2415
rect 4785 -3985 4800 -2415
rect 4500 -4000 4800 -3985
rect 5100 -2415 5400 -2400
rect 5100 -3985 5115 -2415
rect 5385 -3985 5400 -2415
rect 5100 -4000 5400 -3985
rect 5700 -2415 6000 -2400
rect 5700 -3985 5715 -2415
rect 5985 -3985 6000 -2415
rect 5700 -4000 6000 -3985
rect 6300 -2415 6600 -2400
rect 6300 -3985 6315 -2415
rect 6585 -3985 6600 -2415
rect 6300 -4000 6600 -3985
rect 6900 -2415 7200 -2400
rect 6900 -3985 6915 -2415
rect 7185 -3985 7200 -2415
rect 6900 -4000 7200 -3985
rect 7500 -2415 7800 -2400
rect 7500 -3985 7515 -2415
rect 7785 -3985 7800 -2415
rect 7500 -4000 7800 -3985
rect 8100 -2415 8400 -2400
rect 8100 -3985 8115 -2415
rect 8385 -3985 8400 -2415
rect 8100 -4000 8400 -3985
rect 8700 -2415 9000 -2400
rect 8700 -3985 8715 -2415
rect 8985 -3985 9000 -2415
rect 8700 -4000 9000 -3985
rect 9300 -2415 9600 -2400
rect 9300 -3985 9315 -2415
rect 9585 -3985 9600 -2415
rect 9300 -4000 9600 -3985
rect 9900 -2415 10200 -2400
rect 9900 -3985 9915 -2415
rect 10185 -3985 10200 -2415
rect 9900 -4000 10200 -3985
rect 10500 -2415 10800 -2400
rect 10500 -3985 10515 -2415
rect 10785 -3985 10800 -2415
rect 10500 -4000 10800 -3985
rect 11100 -2415 11400 -2400
rect 11100 -3985 11115 -2415
rect 11385 -3985 11400 -2415
rect 11100 -4000 11400 -3985
<< ndiffc >>
rect -285 15 -15 1585
rect 315 15 585 1585
rect 915 15 1185 1585
rect 1515 15 1785 1585
rect 2115 15 2385 1585
rect 2715 15 2985 1585
rect 3315 15 3585 1585
rect 3915 15 4185 1585
rect 4515 15 4785 1585
rect 5115 15 5385 1585
rect 5715 15 5985 1585
rect 6315 15 6585 1585
rect 6915 15 7185 1585
rect 7515 15 7785 1585
rect 8115 15 8385 1585
rect 8715 15 8985 1585
rect 9315 15 9585 1585
rect 9915 15 10185 1585
rect 10515 15 10785 1585
rect 11115 15 11385 1585
rect -285 -1985 -15 -415
rect 315 -1985 585 -415
rect 915 -1985 1185 -415
rect 1515 -1985 1785 -415
rect 2115 -1985 2385 -415
rect 2715 -1985 2985 -415
rect 3315 -1985 3585 -415
rect 3915 -1985 4185 -415
rect 4515 -1985 4785 -415
rect 5115 -1985 5385 -415
rect 5715 -1985 5985 -415
rect 6315 -1985 6585 -415
rect 6915 -1985 7185 -415
rect 7515 -1985 7785 -415
rect 8115 -1985 8385 -415
rect 8715 -1985 8985 -415
rect 9315 -1985 9585 -415
rect 9915 -1985 10185 -415
rect 10515 -1985 10785 -415
rect 11115 -1985 11385 -415
rect -285 -3985 -15 -2415
rect 315 -3985 585 -2415
rect 915 -3985 1185 -2415
rect 1515 -3985 1785 -2415
rect 2115 -3985 2385 -2415
rect 2715 -3985 2985 -2415
rect 3315 -3985 3585 -2415
rect 3915 -3985 4185 -2415
rect 4515 -3985 4785 -2415
rect 5115 -3985 5385 -2415
rect 5715 -3985 5985 -2415
rect 6315 -3985 6585 -2415
rect 6915 -3985 7185 -2415
rect 7515 -3985 7785 -2415
rect 8115 -3985 8385 -2415
rect 8715 -3985 8985 -2415
rect 9315 -3985 9585 -2415
rect 9915 -3985 10185 -2415
rect 10515 -3985 10785 -2415
rect 11115 -3985 11385 -2415
<< psubdiff >>
rect 2225 1665 2275 1680
rect 2225 1645 2240 1665
rect 2260 1645 2275 1665
rect 2825 1665 2875 1680
rect 2225 1630 2275 1645
rect 2825 1645 2840 1665
rect 2860 1645 2875 1665
rect 4625 1665 4675 1680
rect 2825 1630 2875 1645
rect 4625 1645 4640 1665
rect 4660 1645 4675 1665
rect 5225 1665 5275 1680
rect 4625 1630 4675 1645
rect 5225 1645 5240 1665
rect 5260 1645 5275 1665
rect 6425 1665 6475 1680
rect 5225 1630 5275 1645
rect 6425 1645 6440 1665
rect 6460 1645 6475 1665
rect 7625 1665 7675 1680
rect 6425 1630 6475 1645
rect 7625 1645 7640 1665
rect 7660 1645 7675 1665
rect 8825 1665 8875 1680
rect 7625 1630 7675 1645
rect 8825 1645 8840 1665
rect 8860 1645 8875 1665
rect 8825 1630 8875 1645
rect -600 1585 -300 1600
rect -600 15 -585 1585
rect -315 15 -300 1585
rect -600 0 -300 15
rect 11400 1585 11700 1600
rect 11400 15 11415 1585
rect 11685 15 11700 1585
rect 11400 0 11700 15
rect 2225 -155 2275 -140
rect 2225 -175 2240 -155
rect 2260 -175 2275 -155
rect 2225 -190 2275 -175
rect 8225 -205 8275 -190
rect 4025 -235 4075 -220
rect 4025 -255 4040 -235
rect 4060 -255 4075 -235
rect 4025 -270 4075 -255
rect 5825 -235 5875 -220
rect 5825 -255 5840 -235
rect 5860 -255 5875 -235
rect 8225 -225 8240 -205
rect 8260 -225 8275 -205
rect 8225 -240 8275 -225
rect 5825 -270 5875 -255
rect 9425 -235 9475 -220
rect 9425 -255 9440 -235
rect 9460 -255 9475 -235
rect 9425 -270 9475 -255
rect -600 -415 -300 -400
rect -600 -1985 -585 -415
rect -315 -1985 -300 -415
rect -600 -2000 -300 -1985
rect 11400 -415 11700 -400
rect 11400 -1985 11415 -415
rect 11685 -1985 11700 -415
rect 11400 -2000 11700 -1985
rect 1625 -2335 1675 -2320
rect 1625 -2355 1640 -2335
rect 1660 -2355 1675 -2335
rect 1625 -2370 1675 -2355
rect 4025 -2335 4075 -2320
rect 4025 -2355 4040 -2335
rect 4060 -2355 4075 -2335
rect 4025 -2370 4075 -2355
rect 5825 -2330 5875 -2315
rect 5825 -2350 5840 -2330
rect 5860 -2350 5875 -2330
rect 5825 -2365 5875 -2350
rect 7655 -2330 7705 -2315
rect 7655 -2350 7670 -2330
rect 7690 -2350 7705 -2330
rect 7655 -2365 7705 -2350
rect 9425 -2330 9475 -2315
rect 9425 -2350 9440 -2330
rect 9460 -2350 9475 -2330
rect 9425 -2365 9475 -2350
rect -600 -2415 -300 -2400
rect -600 -3985 -585 -2415
rect -315 -3985 -300 -2415
rect -600 -4000 -300 -3985
rect 11400 -2415 11700 -2400
rect 11400 -3985 11415 -2415
rect 11685 -3985 11700 -2415
rect 11400 -4000 11700 -3985
rect 2225 -4045 2275 -4030
rect 2225 -4065 2240 -4045
rect 2260 -4065 2275 -4045
rect 4025 -4045 4075 -4030
rect 2225 -4080 2275 -4065
rect 4025 -4065 4040 -4045
rect 4060 -4065 4075 -4045
rect 5825 -4045 5875 -4030
rect 4025 -4080 4075 -4065
rect 5825 -4065 5840 -4045
rect 5860 -4065 5875 -4045
rect 7625 -4045 7675 -4030
rect 5825 -4080 5875 -4065
rect 7625 -4065 7640 -4045
rect 7660 -4065 7675 -4045
rect 7625 -4080 7675 -4065
rect 9300 -4060 9350 -4055
rect 9300 -4080 9315 -4060
rect 9335 -4080 9350 -4060
rect 9300 -4095 9350 -4080
<< psubdiffcont >>
rect 2240 1645 2260 1665
rect 2840 1645 2860 1665
rect 4640 1645 4660 1665
rect 5240 1645 5260 1665
rect 6440 1645 6460 1665
rect 7640 1645 7660 1665
rect 8840 1645 8860 1665
rect -585 15 -315 1585
rect 11415 15 11685 1585
rect 2240 -175 2260 -155
rect 4040 -255 4060 -235
rect 5840 -255 5860 -235
rect 8240 -225 8260 -205
rect 9440 -255 9460 -235
rect -585 -1985 -315 -415
rect 11415 -1985 11685 -415
rect 1640 -2355 1660 -2335
rect 4040 -2355 4060 -2335
rect 5840 -2350 5860 -2330
rect 7670 -2350 7690 -2330
rect 9440 -2350 9460 -2330
rect -585 -3985 -315 -2415
rect 11415 -3985 11685 -2415
rect 2240 -4065 2260 -4045
rect 4040 -4065 4060 -4045
rect 5840 -4065 5860 -4045
rect 7640 -4065 7660 -4045
rect 9315 -4080 9335 -4060
<< poly >>
rect 9615 1705 9900 1715
rect 9615 1685 9625 1705
rect 9890 1685 9900 1705
rect -295 1645 900 1655
rect -295 1625 -285 1645
rect -15 1625 315 1645
rect 585 1625 900 1645
rect -295 1615 900 1625
rect 0 1600 300 1615
rect 600 1600 900 1615
rect 1200 1640 2225 1655
rect 1200 1600 1500 1640
rect 1800 1600 2100 1640
rect 2275 1640 2825 1655
rect 2875 1640 4625 1655
rect 2400 1600 2700 1615
rect 3000 1600 3300 1640
rect 3600 1600 3900 1615
rect 4200 1600 4500 1640
rect 4675 1640 5225 1655
rect 5275 1640 6425 1655
rect 4800 1600 5100 1615
rect 5400 1600 5700 1640
rect 6475 1640 7625 1655
rect 6000 1600 6300 1615
rect 6600 1600 6900 1640
rect 7675 1640 8825 1655
rect 9615 1655 9900 1685
rect 7200 1600 7500 1615
rect 7800 1600 8100 1640
rect 8875 1640 9900 1655
rect 8400 1600 8700 1615
rect 9000 1600 9300 1640
rect 9600 1600 9900 1640
rect 10200 1645 11395 1655
rect 10200 1625 10515 1645
rect 10785 1625 11115 1645
rect 11385 1625 11395 1645
rect 10200 1615 11395 1625
rect 10200 1600 10500 1615
rect 10800 1600 11100 1615
rect 0 -15 300 0
rect 600 -15 900 0
rect 1200 -15 1500 0
rect 1800 -15 2100 0
rect 2400 -15 2700 0
rect 3000 -15 3300 0
rect 3600 -15 3900 0
rect 4200 -15 4500 0
rect 4800 -15 5100 0
rect 5400 -15 5700 0
rect 6000 -15 6300 0
rect 6600 -15 6900 0
rect 7200 -15 7500 0
rect 7800 -15 8100 0
rect 8400 -15 8700 0
rect 2530 -25 2570 -15
rect 2530 -45 2540 -25
rect 2560 -45 2570 -25
rect 2530 -55 2570 -45
rect 3730 -25 3770 -15
rect 3730 -45 3740 -25
rect 3760 -45 3770 -25
rect 3730 -55 3770 -45
rect 4930 -25 4970 -15
rect 4930 -45 4940 -25
rect 4960 -45 4970 -25
rect 4930 -55 4970 -45
rect 6130 -25 6170 -15
rect 6130 -45 6140 -25
rect 6160 -45 6170 -25
rect 6130 -55 6170 -45
rect 7330 -25 7370 -15
rect 7330 -45 7340 -25
rect 7360 -45 7370 -25
rect 7330 -55 7370 -45
rect 8530 -25 8570 -15
rect 8530 -45 8540 -25
rect 8560 -45 8570 -25
rect 8530 -55 8570 -45
rect 3565 -305 3935 -260
rect 6575 -305 6925 -265
rect 9000 -305 9300 0
rect 9600 -15 9900 0
rect 10200 -15 10500 0
rect 10800 -15 11100 0
rect 1200 -345 3605 -305
rect 3895 -345 6615 -305
rect 6885 -345 9300 -305
rect -295 -355 900 -345
rect -295 -375 -285 -355
rect -15 -375 315 -355
rect 585 -375 900 -355
rect -295 -385 900 -375
rect 0 -400 300 -385
rect 600 -400 900 -385
rect 1200 -400 1500 -345
rect 1800 -400 2100 -345
rect 2400 -400 2700 -345
rect 3000 -400 3300 -345
rect 3730 -355 3770 -345
rect 3730 -375 3740 -355
rect 3760 -375 3770 -355
rect 3730 -385 3770 -375
rect 3600 -400 3900 -385
rect 4200 -400 4500 -345
rect 4800 -400 5100 -345
rect 5400 -400 5700 -345
rect 6000 -400 6300 -345
rect 6730 -355 6770 -345
rect 6730 -375 6740 -355
rect 6760 -375 6770 -355
rect 6730 -385 6770 -375
rect 6600 -400 6900 -385
rect 7200 -400 7500 -345
rect 7800 -400 8100 -345
rect 8400 -400 8700 -345
rect 9000 -400 9300 -345
rect 9905 -355 10195 -345
rect 9905 -370 9915 -355
rect 9600 -375 9915 -370
rect 10185 -370 10195 -355
rect 10505 -355 10795 -345
rect 10505 -370 10515 -355
rect 10185 -375 10515 -370
rect 10785 -370 10795 -355
rect 11105 -355 11395 -345
rect 11105 -370 11115 -355
rect 10785 -375 11115 -370
rect 11385 -375 11395 -355
rect 9600 -385 11395 -375
rect 9600 -400 9900 -385
rect 10200 -400 10500 -385
rect 10800 -400 11100 -385
rect 0 -2015 300 -2000
rect 600 -2015 900 -2000
rect 1200 -2015 1500 -2000
rect 1800 -2015 2100 -2000
rect 2400 -2015 2700 -2000
rect 3000 -2015 3300 -2000
rect 3600 -2015 3900 -2000
rect 4200 -2015 4500 -2000
rect 4800 -2015 5100 -2000
rect 5400 -2015 5700 -2000
rect 6000 -2015 6300 -2000
rect 6600 -2015 6900 -2000
rect 7200 -2015 7500 -2000
rect 7800 -2015 8100 -2000
rect 8400 -2015 8700 -2000
rect 9000 -2015 9300 -2000
rect 9600 -2015 9900 -2000
rect 10200 -2015 10500 -2000
rect 10800 -2015 11100 -2000
rect 1735 -2025 1775 -2015
rect 1735 -2045 1745 -2025
rect 1765 -2045 1775 -2025
rect 1735 -2345 1775 -2045
rect 4630 -2025 4670 -2015
rect 4630 -2045 4640 -2025
rect 4660 -2045 4670 -2025
rect 1735 -2365 1745 -2345
rect 1765 -2365 1775 -2345
rect 1735 -2375 1775 -2365
rect 4630 -2355 4670 -2045
rect 7525 -2025 7565 -2015
rect 7525 -2045 7535 -2025
rect 7555 -2045 7565 -2025
rect 7525 -2285 7565 -2045
rect 7525 -2305 7535 -2285
rect 7555 -2305 7565 -2285
rect 7525 -2315 7565 -2305
rect 8725 -2025 8765 -2015
rect 8725 -2045 8735 -2025
rect 8755 -2045 8765 -2025
rect 4630 -2375 4640 -2355
rect 4660 -2375 4670 -2355
rect 8725 -2350 8765 -2045
rect 4630 -2385 4670 -2375
rect 8725 -2370 8735 -2350
rect 8755 -2370 8765 -2350
rect 8725 -2380 8765 -2370
rect 0 -2400 300 -2385
rect 600 -2400 900 -2385
rect 1200 -2400 1500 -2385
rect 1800 -2400 2100 -2385
rect 2400 -2400 2700 -2385
rect 3000 -2400 3300 -2385
rect 3600 -2400 3900 -2385
rect 4200 -2400 4500 -2385
rect 4800 -2400 5100 -2385
rect 5400 -2400 5700 -2385
rect 6000 -2400 6300 -2385
rect 6600 -2400 6900 -2385
rect 7200 -2400 7500 -2385
rect 7800 -2400 8100 -2385
rect 8400 -2400 8700 -2385
rect 9000 -2400 9300 -2385
rect 9600 -2400 9900 -2385
rect 10200 -2400 10500 -2385
rect 10800 -2400 11100 -2385
rect 0 -4015 300 -4000
rect 600 -4015 900 -4000
rect 1200 -4015 1500 -4000
rect 1800 -4015 2100 -4000
rect 2400 -4015 2700 -4000
rect -295 -4025 2100 -4015
rect -295 -4045 -285 -4025
rect -15 -4045 315 -4025
rect 585 -4045 915 -4025
rect 1185 -4045 1515 -4025
rect 1785 -4045 2100 -4025
rect 3000 -4025 3300 -4000
rect -295 -4055 2100 -4045
rect 3000 -4045 3010 -4025
rect 3290 -4045 3300 -4025
rect 3000 -4055 3300 -4045
rect 3600 -4025 3900 -4000
rect 3600 -4045 3740 -4025
rect 3760 -4045 3900 -4025
rect 4200 -4025 4500 -4000
rect 3600 -4055 3900 -4045
rect 4200 -4045 4210 -4025
rect 4490 -4045 4500 -4025
rect 4200 -4055 4500 -4045
rect 4800 -4025 5100 -4000
rect 4800 -4045 4810 -4025
rect 5090 -4045 5100 -4025
rect 4800 -4055 5100 -4045
rect 5400 -4025 5700 -4000
rect 5400 -4045 5410 -4025
rect 5690 -4045 5700 -4025
rect 6000 -4025 6300 -4000
rect 5400 -4055 5700 -4045
rect 6000 -4045 6010 -4025
rect 6285 -4045 6300 -4025
rect 6000 -4055 6300 -4045
rect 6600 -4025 6900 -4000
rect 6600 -4045 6605 -4025
rect 6890 -4045 6900 -4025
rect 6600 -4055 6900 -4045
rect 7200 -4025 7500 -4000
rect 7200 -4045 7210 -4025
rect 7490 -4045 7500 -4025
rect 7800 -4025 8100 -4000
rect 7200 -4055 7500 -4045
rect 7800 -4045 7810 -4025
rect 8090 -4045 8100 -4025
rect 7800 -4055 8100 -4045
rect 8400 -4015 8700 -4000
rect 9000 -4015 9300 -4000
rect 9600 -4015 9900 -4000
rect 10200 -4015 10500 -4000
rect 10800 -4015 11100 -4000
rect 8400 -4025 11395 -4015
rect 8400 -4045 8715 -4025
rect 8985 -4045 9385 -4025
rect 9585 -4045 9915 -4025
rect 10185 -4045 10515 -4025
rect 10785 -4045 11115 -4025
rect 11385 -4045 11395 -4025
rect 8400 -4055 11395 -4045
<< polycont >>
rect 9625 1685 9890 1705
rect -285 1625 -15 1645
rect 315 1625 585 1645
rect 10515 1625 10785 1645
rect 11115 1625 11385 1645
rect 2540 -45 2560 -25
rect 3740 -45 3760 -25
rect 4940 -45 4960 -25
rect 6140 -45 6160 -25
rect 7340 -45 7360 -25
rect 8540 -45 8560 -25
rect -285 -375 -15 -355
rect 315 -375 585 -355
rect 3740 -375 3760 -355
rect 6740 -375 6760 -355
rect 9915 -375 10185 -355
rect 10515 -375 10785 -355
rect 11115 -375 11385 -355
rect 1745 -2045 1765 -2025
rect 4640 -2045 4660 -2025
rect 1745 -2365 1765 -2345
rect 7535 -2045 7555 -2025
rect 7535 -2305 7555 -2285
rect 8735 -2045 8755 -2025
rect 4640 -2375 4660 -2355
rect 8735 -2370 8755 -2350
rect -285 -4045 -15 -4025
rect 315 -4045 585 -4025
rect 915 -4045 1185 -4025
rect 1515 -4045 1785 -4025
rect 3010 -4045 3290 -4025
rect 3740 -4045 3760 -4025
rect 4210 -4045 4490 -4025
rect 4810 -4045 5090 -4025
rect 5410 -4045 5690 -4025
rect 6010 -4045 6285 -4025
rect 6605 -4045 6890 -4025
rect 7210 -4045 7490 -4025
rect 7810 -4045 8090 -4025
rect 8715 -4045 8985 -4025
rect 9385 -4045 9585 -4025
rect 9915 -4045 10185 -4025
rect 10515 -4045 10785 -4025
rect 11115 -4045 11385 -4025
<< locali >>
rect 9305 1740 11700 1780
rect 2230 1665 2270 1675
rect -295 1645 -5 1655
rect -295 1625 -285 1645
rect -15 1625 -5 1645
rect -295 1595 -5 1625
rect -595 1585 -5 1595
rect -595 15 -585 1585
rect -315 15 -285 1585
rect -15 15 -5 1585
rect -595 5 -5 15
rect 305 1645 595 1655
rect 305 1625 315 1645
rect 585 1625 595 1645
rect 2230 1645 2240 1665
rect 2260 1645 2270 1665
rect 2230 1635 2270 1645
rect 2830 1665 2870 1675
rect 2830 1645 2840 1665
rect 2860 1645 2870 1665
rect 2830 1635 2870 1645
rect 4630 1665 4670 1675
rect 4630 1645 4640 1665
rect 4660 1645 4670 1665
rect 4630 1635 4670 1645
rect 5230 1665 5270 1675
rect 5230 1645 5240 1665
rect 5260 1645 5270 1665
rect 5230 1635 5270 1645
rect 6430 1665 6470 1675
rect 6430 1645 6440 1665
rect 6460 1645 6470 1665
rect 6430 1635 6470 1645
rect 7630 1665 7670 1675
rect 7630 1645 7640 1665
rect 7660 1645 7670 1665
rect 7630 1635 7670 1645
rect 8830 1665 8870 1675
rect 8830 1645 8840 1665
rect 8860 1645 8870 1665
rect 8830 1635 8870 1645
rect 305 1585 595 1625
rect 305 15 315 1585
rect 585 15 595 1585
rect 305 5 595 15
rect 905 1585 1195 1595
rect 905 15 915 1585
rect 1185 15 1195 1585
rect 905 -20 1195 15
rect 1505 1585 1795 1595
rect 1505 15 1515 1585
rect 1785 15 1795 1585
rect 1505 5 1795 15
rect 2105 1585 2400 1595
rect 2105 15 2115 1585
rect 2385 15 2400 1585
rect 2105 5 2400 15
rect 2705 1585 2995 1595
rect 2705 15 2715 1585
rect 2985 15 2995 1585
rect 2105 -20 2395 5
rect 905 -60 2395 -20
rect 2530 -25 2570 -15
rect 2530 -45 2540 -25
rect 2560 -45 2570 -25
rect 2705 -40 2995 15
rect 3305 1585 3595 1595
rect 3305 15 3315 1585
rect 3585 15 3595 1585
rect 3305 5 3595 15
rect 3905 1585 4195 1595
rect 3905 15 3915 1585
rect 4185 15 4195 1585
rect 3905 5 4195 15
rect 4505 1585 4795 1595
rect 4505 15 4515 1585
rect 4785 15 4795 1585
rect 3730 -25 3770 -15
rect 2530 -55 2570 -45
rect -295 -355 -5 -345
rect -295 -375 -285 -355
rect -15 -375 -5 -355
rect -295 -405 -5 -375
rect -595 -415 -5 -405
rect -595 -1985 -585 -415
rect -315 -1985 -285 -415
rect -15 -1985 -5 -415
rect -595 -1995 -5 -1985
rect 305 -355 595 -345
rect 305 -375 315 -355
rect 585 -375 595 -355
rect 305 -415 595 -375
rect 305 -1985 315 -415
rect 585 -1985 595 -415
rect 305 -1995 595 -1985
rect 905 -415 1195 -405
rect 905 -1985 915 -415
rect 1185 -1985 1195 -415
rect 905 -2080 1195 -1985
rect 1505 -415 1795 -60
rect 2230 -155 2270 -145
rect 2230 -175 2240 -155
rect 2260 -175 2270 -155
rect 2230 -185 2270 -175
rect 2820 -255 2860 -40
rect 3730 -45 3740 -25
rect 3760 -45 3770 -25
rect 3730 -55 3770 -45
rect 1505 -1985 1515 -415
rect 1785 -1985 1795 -415
rect 1505 -2015 1795 -1985
rect 2105 -295 2860 -255
rect 4030 -235 4070 -220
rect 4030 -255 4040 -235
rect 4060 -255 4070 -235
rect 4030 -265 4070 -255
rect 2105 -405 2395 -295
rect 3580 -320 3920 -280
rect 4505 -320 4795 15
rect 5105 1585 5395 1595
rect 5105 15 5115 1585
rect 5385 15 5395 1585
rect 4930 -25 4970 -15
rect 4930 -45 4940 -25
rect 4960 -45 4970 -25
rect 4930 -55 4970 -45
rect 2705 -360 3620 -320
rect 3730 -355 3770 -345
rect 2105 -415 2400 -405
rect 2105 -1985 2115 -415
rect 2385 -1985 2400 -415
rect 2105 -1995 2400 -1985
rect 2705 -415 2995 -360
rect 3730 -375 3740 -355
rect 3760 -375 3770 -355
rect 3880 -360 4795 -320
rect 3730 -385 3770 -375
rect 2705 -1985 2715 -415
rect 2985 -1985 2995 -415
rect 2705 -1995 2995 -1985
rect 3305 -415 3595 -405
rect 3305 -1985 3315 -415
rect 3585 -1985 3595 -415
rect 1735 -2025 1775 -2015
rect 1735 -2045 1745 -2025
rect 1765 -2045 1775 -2025
rect 1735 -2055 1775 -2045
rect 2105 -2080 2395 -1995
rect 3305 -2080 3595 -1985
rect 905 -2120 3595 -2080
rect 3905 -415 4195 -405
rect 3905 -1985 3915 -415
rect 4185 -1985 4195 -415
rect 3905 -2080 4195 -1985
rect 4505 -415 4795 -360
rect 4505 -1985 4515 -415
rect 4785 -1985 4795 -415
rect 4505 -2015 4795 -1985
rect 5105 -320 5395 15
rect 5705 1585 5995 1595
rect 5705 15 5715 1585
rect 5985 15 5995 1585
rect 5705 5 5995 15
rect 6305 1585 6595 1595
rect 6305 15 6315 1585
rect 6585 15 6595 1585
rect 6130 -25 6170 -15
rect 6130 -45 6140 -25
rect 6160 -45 6170 -25
rect 6130 -55 6170 -45
rect 5830 -235 5870 -225
rect 5830 -255 5840 -235
rect 5860 -255 5870 -235
rect 5830 -265 5870 -255
rect 6305 -260 6595 15
rect 6905 1585 7195 1595
rect 6905 15 6915 1585
rect 7185 15 7195 1585
rect 6905 5 7195 15
rect 7505 1585 7795 1595
rect 7505 15 7515 1585
rect 7785 15 7795 1585
rect 7330 -25 7370 -15
rect 7330 -45 7340 -25
rect 7360 -45 7370 -25
rect 7330 -55 7370 -45
rect 7505 -260 7795 15
rect 8105 1585 8395 1595
rect 8105 15 8115 1585
rect 8385 15 8395 1585
rect 8105 5 8395 15
rect 8705 1585 8995 1595
rect 8705 15 8715 1585
rect 8985 15 8995 1585
rect 8530 -25 8570 -15
rect 8530 -45 8540 -25
rect 8560 -45 8570 -25
rect 8530 -55 8570 -45
rect 8705 -20 8995 15
rect 9305 1585 9595 1740
rect 9615 1705 11700 1715
rect 9615 1685 9625 1705
rect 9890 1685 11700 1705
rect 9615 1675 11700 1685
rect 10505 1645 10795 1655
rect 10505 1625 10515 1645
rect 10785 1625 10795 1645
rect 9305 15 9315 1585
rect 9585 15 9595 1585
rect 9305 5 9595 15
rect 9905 1585 10195 1595
rect 9905 15 9915 1585
rect 10185 15 10195 1585
rect 9905 -20 10195 15
rect 10505 1585 10795 1625
rect 10505 15 10515 1585
rect 10785 15 10795 1585
rect 10505 5 10795 15
rect 11105 1645 11395 1655
rect 11105 1625 11115 1645
rect 11385 1625 11395 1645
rect 11105 1595 11395 1625
rect 11105 1585 11695 1595
rect 11105 15 11115 1585
rect 11385 15 11415 1585
rect 11685 15 11695 1585
rect 11105 5 11695 15
rect 8705 -60 10195 -20
rect 8230 -205 8270 -195
rect 8230 -225 8240 -205
rect 8260 -225 8270 -205
rect 8230 -235 8270 -225
rect 6305 -300 6920 -260
rect 7505 -300 8395 -260
rect 6880 -320 6920 -300
rect 5105 -360 6595 -320
rect 5105 -415 5395 -360
rect 5105 -1985 5115 -415
rect 5385 -1985 5395 -415
rect 4630 -2025 4670 -2015
rect 4630 -2045 4640 -2025
rect 4660 -2045 4670 -2025
rect 4630 -2055 4670 -2045
rect 5105 -2080 5395 -1985
rect 5705 -415 5995 -405
rect 5705 -1985 5715 -415
rect 5985 -1985 5995 -415
rect 5705 -2015 5995 -1985
rect 6305 -415 6595 -360
rect 6730 -355 6770 -345
rect 6730 -375 6740 -355
rect 6760 -375 6770 -355
rect 6880 -360 7795 -320
rect 6730 -385 6770 -375
rect 6305 -1985 6315 -415
rect 6585 -1985 6595 -415
rect 6305 -1995 6595 -1985
rect 6905 -415 7195 -405
rect 6905 -1985 6915 -415
rect 7185 -1985 7195 -415
rect 3905 -2120 5395 -2080
rect 1630 -2335 1670 -2325
rect 1630 -2355 1640 -2335
rect 1660 -2355 1670 -2335
rect 1630 -2405 1670 -2355
rect 1735 -2345 2995 -2335
rect 1735 -2365 1745 -2345
rect 1765 -2365 2995 -2345
rect 1735 -2375 2995 -2365
rect -595 -2415 -5 -2405
rect -595 -3985 -585 -2415
rect -315 -3985 -285 -2415
rect -15 -3985 -5 -2415
rect -595 -3995 -5 -3985
rect -295 -4025 -5 -3995
rect -295 -4045 -285 -4025
rect -15 -4045 -5 -4025
rect -295 -4055 -5 -4045
rect 305 -2415 595 -2405
rect 305 -3985 315 -2415
rect 585 -3985 595 -2415
rect 305 -4025 595 -3985
rect 305 -4045 315 -4025
rect 585 -4045 595 -4025
rect 305 -4055 595 -4045
rect 905 -2415 1195 -2405
rect 905 -3985 915 -2415
rect 1185 -3985 1195 -2415
rect 905 -4025 1195 -3985
rect 905 -4045 915 -4025
rect 1185 -4045 1195 -4025
rect 905 -4055 1195 -4045
rect 1505 -2415 1795 -2405
rect 1505 -3985 1515 -2415
rect 1785 -3985 1795 -2415
rect 1505 -4025 1795 -3985
rect 2105 -2415 2400 -2405
rect 2105 -3985 2115 -2415
rect 2385 -3985 2400 -2415
rect 2105 -3995 2400 -3985
rect 2705 -2415 2995 -2375
rect 2705 -3985 2715 -2415
rect 2985 -3985 2995 -2415
rect 2705 -3995 2995 -3985
rect 3305 -2415 3595 -2120
rect 4030 -2335 4070 -2325
rect 4030 -2355 4040 -2335
rect 4060 -2355 4070 -2335
rect 4030 -2405 4070 -2355
rect 4630 -2355 4670 -2345
rect 4630 -2375 4640 -2355
rect 4660 -2375 4670 -2355
rect 4630 -2385 4670 -2375
rect 3305 -3985 3315 -2415
rect 3585 -3985 3595 -2415
rect 3305 -3995 3595 -3985
rect 3905 -2415 4195 -2405
rect 3905 -3985 3915 -2415
rect 4185 -3985 4195 -2415
rect 3905 -3995 4195 -3985
rect 4505 -2415 4795 -2385
rect 4505 -3985 4515 -2415
rect 4785 -3985 4795 -2415
rect 4505 -3995 4795 -3985
rect 5105 -2415 5395 -2120
rect 5955 -2275 5995 -2015
rect 6905 -2080 7195 -1985
rect 7505 -415 7795 -360
rect 7505 -1985 7515 -415
rect 7785 -1985 7795 -415
rect 7505 -2015 7795 -1985
rect 8105 -415 8395 -300
rect 8105 -1985 8115 -415
rect 8385 -1985 8395 -415
rect 7525 -2025 7565 -2015
rect 7525 -2045 7535 -2025
rect 7555 -2045 7565 -2025
rect 7525 -2055 7565 -2045
rect 8105 -2080 8395 -1985
rect 8705 -415 8995 -60
rect 9430 -235 9470 -225
rect 9430 -255 9440 -235
rect 9460 -255 9470 -235
rect 9430 -265 9470 -255
rect 9905 -355 10195 -345
rect 9905 -375 9915 -355
rect 10185 -375 10195 -355
rect 8705 -1985 8715 -415
rect 8985 -1985 8995 -415
rect 8705 -2015 8995 -1985
rect 9305 -415 9595 -405
rect 9305 -1985 9315 -415
rect 9585 -1985 9595 -415
rect 8725 -2025 8765 -2015
rect 8725 -2045 8735 -2025
rect 8755 -2045 8765 -2025
rect 8725 -2055 8765 -2045
rect 9305 -2080 9595 -1985
rect 9905 -415 10195 -375
rect 9905 -1985 9915 -415
rect 10185 -1985 10195 -415
rect 9905 -1995 10195 -1985
rect 10505 -355 10795 -345
rect 10505 -375 10515 -355
rect 10785 -375 10795 -355
rect 10505 -415 10795 -375
rect 10505 -1985 10515 -415
rect 10785 -1985 10795 -415
rect 10505 -1995 10795 -1985
rect 11105 -355 11395 -345
rect 11105 -375 11115 -355
rect 11385 -375 11395 -355
rect 11105 -405 11395 -375
rect 11105 -415 11695 -405
rect 11105 -1985 11115 -415
rect 11385 -1985 11415 -415
rect 11685 -1985 11695 -415
rect 11105 -1995 11695 -1985
rect 6905 -2120 9595 -2080
rect 5955 -2285 7565 -2275
rect 5955 -2305 7535 -2285
rect 7555 -2305 7565 -2285
rect 5955 -2315 7565 -2305
rect 5830 -2330 5870 -2320
rect 5830 -2350 5840 -2330
rect 5860 -2350 5870 -2330
rect 5830 -2405 5870 -2350
rect 5105 -3985 5115 -2415
rect 5385 -3985 5395 -2415
rect 5105 -3995 5395 -3985
rect 5705 -2415 5995 -2405
rect 5705 -3985 5715 -2415
rect 5985 -3985 5995 -2415
rect 5705 -3995 5995 -3985
rect 6305 -2415 6595 -2315
rect 7585 -2340 7625 -2120
rect 6305 -3985 6315 -2415
rect 6585 -3985 6595 -2415
rect 6305 -3995 6595 -3985
rect 6905 -2380 7625 -2340
rect 7660 -2330 7700 -2320
rect 7660 -2350 7670 -2330
rect 7690 -2350 7700 -2330
rect 9430 -2330 9470 -2320
rect 6905 -2415 7195 -2380
rect 7660 -2405 7700 -2350
rect 8725 -2350 8765 -2340
rect 8725 -2360 8735 -2350
rect 8105 -2370 8735 -2360
rect 8755 -2370 8765 -2350
rect 8105 -2380 8765 -2370
rect 9430 -2350 9440 -2330
rect 9460 -2350 9470 -2330
rect 6905 -3985 6915 -2415
rect 7185 -3985 7195 -2415
rect 6905 -3995 7195 -3985
rect 7505 -2415 7795 -2405
rect 7505 -3985 7515 -2415
rect 7785 -3985 7795 -2415
rect 7505 -3995 7795 -3985
rect 8105 -2415 8395 -2380
rect 9430 -2405 9470 -2350
rect 8105 -3985 8115 -2415
rect 8385 -3985 8395 -2415
rect 8105 -3995 8395 -3985
rect 8705 -2415 8995 -2405
rect 8705 -3985 8715 -2415
rect 8985 -3985 8995 -2415
rect 1505 -4045 1515 -4025
rect 1785 -4045 1795 -4025
rect 1505 -4055 1795 -4045
rect 2230 -4045 2270 -3995
rect 2230 -4065 2240 -4045
rect 2260 -4065 2270 -4045
rect 3000 -4025 3300 -4015
rect 3000 -4045 3010 -4025
rect 3290 -4045 3300 -4025
rect 3000 -4055 3300 -4045
rect 3730 -4025 3770 -4015
rect 3730 -4045 3740 -4025
rect 3760 -4045 3770 -4025
rect 3730 -4055 3770 -4045
rect 4030 -4045 4070 -3995
rect 2230 -4075 2270 -4065
rect 4030 -4065 4040 -4045
rect 4060 -4065 4070 -4045
rect 4200 -4025 4500 -4015
rect 4200 -4045 4210 -4025
rect 4490 -4045 4500 -4025
rect 4200 -4055 4500 -4045
rect 4800 -4025 5100 -4015
rect 4800 -4045 4810 -4025
rect 5090 -4045 5100 -4025
rect 4800 -4055 5100 -4045
rect 5400 -4025 5700 -4015
rect 5400 -4045 5410 -4025
rect 5690 -4045 5700 -4025
rect 5400 -4055 5700 -4045
rect 5830 -4045 5870 -3995
rect 4030 -4075 4070 -4065
rect 5830 -4065 5840 -4045
rect 5860 -4065 5870 -4045
rect 6000 -4025 6295 -4015
rect 6000 -4045 6010 -4025
rect 6285 -4045 6295 -4025
rect 6000 -4055 6295 -4045
rect 6600 -4025 6900 -4015
rect 6600 -4045 6605 -4025
rect 6890 -4045 6900 -4025
rect 6600 -4055 6900 -4045
rect 7200 -4025 7500 -4015
rect 7200 -4045 7210 -4025
rect 7490 -4045 7500 -4025
rect 7200 -4055 7500 -4045
rect 7630 -4045 7670 -3995
rect 5830 -4075 5870 -4065
rect 7630 -4065 7640 -4045
rect 7660 -4065 7670 -4045
rect 7800 -4025 8100 -4015
rect 7800 -4045 7810 -4025
rect 8090 -4045 8100 -4025
rect 7800 -4055 8100 -4045
rect 8705 -4025 8995 -3985
rect 8705 -4045 8715 -4025
rect 8985 -4045 8995 -4025
rect 8705 -4055 8995 -4045
rect 9305 -2415 9595 -2405
rect 9305 -3985 9315 -2415
rect 9585 -3985 9595 -2415
rect 9305 -4015 9595 -3985
rect 7630 -4075 7670 -4065
rect 9305 -4060 9345 -4015
rect 9375 -4025 9595 -4015
rect 9375 -4045 9385 -4025
rect 9585 -4045 9595 -4025
rect 9375 -4055 9595 -4045
rect 9905 -2415 10195 -2405
rect 9905 -3985 9915 -2415
rect 10185 -3985 10195 -2415
rect 9905 -4025 10195 -3985
rect 9905 -4045 9915 -4025
rect 10185 -4045 10195 -4025
rect 9905 -4055 10195 -4045
rect 10505 -2415 10795 -2405
rect 10505 -3985 10515 -2415
rect 10785 -3985 10795 -2415
rect 10505 -4025 10795 -3985
rect 10505 -4045 10515 -4025
rect 10785 -4045 10795 -4025
rect 10505 -4055 10795 -4045
rect 11105 -2415 11695 -2405
rect 11105 -3985 11115 -2415
rect 11385 -3985 11415 -2415
rect 11685 -3985 11695 -2415
rect 11105 -3995 11695 -3985
rect 11105 -4025 11395 -3995
rect 11105 -4045 11115 -4025
rect 11385 -4045 11395 -4025
rect 11105 -4055 11395 -4045
rect 9305 -4080 9315 -4060
rect 9335 -4080 9345 -4060
rect 9305 -4090 9345 -4080
<< viali >>
rect -585 15 -315 1585
rect -285 15 -15 1585
rect 2240 1645 2260 1665
rect 2840 1645 2860 1665
rect 4640 1645 4660 1665
rect 5240 1645 5260 1665
rect 6440 1645 6460 1665
rect 7640 1645 7660 1665
rect 8840 1645 8860 1665
rect 315 15 585 1585
rect 1515 15 1785 1585
rect 2540 -45 2560 -25
rect 3315 15 3585 1585
rect 3915 15 4185 1585
rect -585 -1985 -315 -415
rect -285 -1985 -15 -415
rect 315 -1985 585 -415
rect 2240 -175 2260 -155
rect 3740 -45 3760 -25
rect 4040 -255 4060 -235
rect 4940 -45 4960 -25
rect 3740 -375 3760 -355
rect 5715 15 5985 1585
rect 6140 -45 6160 -25
rect 5840 -255 5860 -235
rect 6915 15 7185 1585
rect 7340 -45 7360 -25
rect 8115 15 8385 1585
rect 8540 -45 8560 -25
rect 10515 15 10785 1585
rect 11115 15 11385 1585
rect 11415 15 11685 1585
rect 8240 -225 8260 -205
rect 6740 -375 6760 -355
rect -585 -3985 -315 -2415
rect -285 -3985 -15 -2415
rect 315 -3985 585 -2415
rect 915 -3985 1185 -2415
rect 1515 -3985 1785 -2415
rect 2115 -3985 2385 -2415
rect 3915 -3985 4185 -2415
rect 9440 -255 9460 -235
rect 9915 -1985 10185 -415
rect 10515 -1985 10785 -415
rect 11115 -1985 11385 -415
rect 11415 -1985 11685 -415
rect 5715 -3985 5985 -2415
rect 7515 -3985 7785 -2415
rect 8715 -3985 8985 -2415
rect 3010 -4045 3290 -4025
rect 3740 -4045 3760 -4025
rect 4210 -4045 4490 -4025
rect 4810 -4045 5090 -4025
rect 5410 -4045 5690 -4025
rect 6010 -4045 6285 -4025
rect 6605 -4045 6890 -4025
rect 7210 -4045 7490 -4025
rect 7810 -4045 8090 -4025
rect 9315 -3985 9585 -2415
rect 9915 -3985 10185 -2415
rect 10515 -3985 10785 -2415
rect 11115 -3985 11385 -2415
rect 11415 -3985 11685 -2415
<< metal1 >>
rect -600 1815 11700 3405
rect -600 1585 595 1595
rect -600 15 -585 1585
rect -315 15 -285 1585
rect -15 15 315 1585
rect 585 15 595 1585
rect -600 -400 595 15
rect 1505 1585 1795 1815
rect 1505 15 1515 1585
rect 1785 15 1795 1585
rect 1505 5 1795 15
rect 2105 1665 2395 1690
rect 2105 1645 2240 1665
rect 2260 1645 2395 1665
rect 2105 -155 2395 1645
rect 2705 1665 2995 1690
rect 2705 1645 2840 1665
rect 2860 1645 2995 1665
rect 2105 -175 2240 -155
rect 2260 -175 2395 -155
rect 2105 -400 2395 -175
rect 2530 -25 2570 -15
rect 2530 -45 2540 -25
rect 2560 -45 2570 -25
rect 2530 -400 2570 -45
rect 2705 -400 2995 1645
rect 3305 1585 3595 1815
rect 3305 15 3315 1585
rect 3585 15 3595 1585
rect 3305 5 3595 15
rect 3905 1585 4195 1815
rect 4505 1665 4795 1730
rect 4505 1645 4640 1665
rect 4660 1645 4795 1665
rect 4505 1600 4795 1645
rect 5105 1665 5395 1690
rect 5105 1645 5240 1665
rect 5260 1645 5395 1665
rect 5105 1600 5395 1645
rect 3905 15 3915 1585
rect 4185 15 4195 1585
rect 5705 1585 5995 1815
rect 3905 5 4195 15
rect 3730 -25 3770 -15
rect 3730 -45 3740 -25
rect 3760 -45 3770 -25
rect 3730 -305 3770 -45
rect 3905 -235 4195 -210
rect 3905 -255 4040 -235
rect 4060 -255 4195 -235
rect 3730 -355 3770 -320
rect 3730 -375 3740 -355
rect 3760 -375 3770 -355
rect 3730 -400 3770 -375
rect 3905 -400 4195 -255
rect 4505 -400 4795 1565
rect 4930 -25 4970 -15
rect 4930 -45 4940 -25
rect 4960 -45 4970 -25
rect 4930 -400 4970 -45
rect 5105 -320 5395 1570
rect 5705 15 5715 1585
rect 5985 15 5995 1585
rect 5705 5 5995 15
rect 6305 1665 6595 1690
rect 6305 1645 6440 1665
rect 6460 1645 6595 1665
rect 6130 -25 6170 -15
rect 6130 -45 6140 -25
rect 6160 -45 6170 -25
rect 5705 -235 5995 -210
rect 5705 -255 5840 -235
rect 5860 -255 5995 -235
rect 5705 -320 5995 -255
rect 6130 -320 6170 -45
rect 6305 -320 6595 1645
rect 6905 1585 7195 1815
rect 6905 15 6915 1585
rect 7185 15 7195 1585
rect 6905 5 7195 15
rect 7505 1665 7795 1690
rect 7505 1645 7640 1665
rect 7660 1645 7795 1665
rect 5105 -340 6595 -320
rect 5105 -400 5395 -340
rect 5705 -400 5995 -340
rect 6130 -400 6170 -340
rect 6305 -400 6595 -340
rect 7330 -25 7370 -15
rect 7330 -45 7340 -25
rect 7360 -45 7370 -25
rect 6730 -355 6770 -345
rect 6730 -375 6740 -355
rect 6760 -375 6770 -355
rect 6730 -400 6770 -375
rect 7330 -400 7370 -45
rect 7505 -320 7795 1645
rect 8105 1585 8395 1815
rect 8105 15 8115 1585
rect 8385 15 8395 1585
rect 8105 5 8395 15
rect 8705 1665 8995 1690
rect 8705 1645 8840 1665
rect 8860 1645 8995 1665
rect 8530 -25 8570 -15
rect 8530 -45 8540 -25
rect 8560 -45 8570 -25
rect 7485 -340 7795 -320
rect 7505 -400 7795 -340
rect 8105 -205 8395 -170
rect 8105 -225 8240 -205
rect 8260 -225 8395 -205
rect 8105 -400 8395 -225
rect 8530 -400 8570 -45
rect 8705 -400 8995 1645
rect 10505 1585 11695 1595
rect 10505 15 10515 1585
rect 10785 15 11115 1585
rect 11385 15 11415 1585
rect 11685 15 11695 1585
rect 9305 -235 9595 -175
rect 9305 -255 9440 -235
rect 9460 -255 9595 -235
rect 9305 -400 9595 -255
rect 10505 -400 11695 15
rect -600 -415 11700 -400
rect -600 -1985 -585 -415
rect -315 -1985 -285 -415
rect -15 -1985 315 -415
rect 585 -1985 9915 -415
rect 10185 -1985 10515 -415
rect 10785 -1985 11115 -415
rect 11385 -1985 11415 -415
rect 11685 -1985 11700 -415
rect -600 -2415 11700 -1985
rect -600 -3985 -585 -2415
rect -315 -3985 -285 -2415
rect -15 -3985 315 -2415
rect 585 -3985 915 -2415
rect 1185 -3985 1515 -2415
rect 1785 -3985 2115 -2415
rect 2385 -3985 3915 -2415
rect 4185 -3985 5715 -2415
rect 5985 -3985 7515 -2415
rect 7785 -3985 8715 -2415
rect 8985 -3985 9315 -2415
rect 9585 -3985 9915 -2415
rect 10185 -3985 10515 -2415
rect 10785 -3985 11115 -2415
rect 11385 -3985 11415 -2415
rect 11685 -3985 11700 -2415
rect -600 -3995 11700 -3985
rect 3000 -4025 3300 -3995
rect 3000 -4045 3010 -4025
rect 3290 -4045 3300 -4025
rect 3000 -4055 3300 -4045
rect 3600 -4025 3900 -3995
rect 3600 -4045 3740 -4025
rect 3760 -4045 3900 -4025
rect 3600 -4055 3900 -4045
rect 4200 -4025 4500 -3995
rect 4200 -4045 4210 -4025
rect 4490 -4045 4500 -4025
rect 4200 -4055 4500 -4045
rect 4800 -4025 5100 -3995
rect 4800 -4045 4810 -4025
rect 5090 -4045 5100 -4025
rect 4800 -4055 5100 -4045
rect 5400 -4025 5700 -3995
rect 5400 -4045 5410 -4025
rect 5690 -4045 5700 -4025
rect 5400 -4055 5700 -4045
rect 6000 -4025 6300 -3995
rect 6000 -4045 6010 -4025
rect 6285 -4045 6300 -4025
rect 6000 -4055 6300 -4045
rect 6600 -4025 6900 -3995
rect 6600 -4045 6605 -4025
rect 6890 -4045 6900 -4025
rect 6600 -4055 6900 -4045
rect 7200 -4025 7500 -3995
rect 7200 -4045 7210 -4025
rect 7490 -4045 7500 -4025
rect 7200 -4055 7500 -4045
rect 7800 -4025 8100 -3995
rect 7800 -4045 7810 -4025
rect 8090 -4045 8100 -4025
rect 7800 -4055 8100 -4045
<< end >>
