magic
tech sky130A
timestamp 1617312088
<< nmos >>
rect 0 5 400 1605
rect 800 5 1200 1605
rect 1600 5 2000 1605
rect 2400 5 2800 1605
rect 3200 5 3600 1605
rect 4000 5 4400 1605
rect 4800 5 5200 1605
rect 5600 5 6000 1605
rect 6400 5 6800 1605
rect 7200 5 7600 1605
rect 8000 5 8400 1605
rect 8800 5 9200 1605
rect 9600 5 10000 1605
rect 10400 5 10800 1605
rect 12000 5 12400 1605
rect 12800 5 13200 1605
rect 13600 5 14000 1605
rect 14400 5 14800 1605
rect 15200 5 15600 1605
rect 16000 5 16400 1605
rect 16800 5 17200 1605
rect 17600 5 18000 1605
rect 18400 5 18800 1605
rect 19200 5 19600 1605
rect 20000 5 20400 1605
rect 0 -2395 400 -795
rect 800 -2395 1200 -795
rect 1600 -2395 2000 -795
rect 2400 -2395 2800 -795
rect 3200 -2395 3600 -795
rect 4000 -2395 4400 -795
rect 4800 -2395 5200 -795
rect 5600 -2395 6000 -795
rect 6400 -2395 6800 -795
rect 7200 -2395 7600 -795
rect 8000 -2395 8400 -795
rect 8800 -2395 9200 -795
rect 9600 -2395 10000 -795
rect 10400 -2395 10800 -795
rect 0 -4795 400 -3195
rect 800 -4795 1200 -3195
rect 1600 -4795 2000 -3195
rect 2400 -4795 2800 -3195
rect 3200 -4795 3600 -3195
rect 4000 -4795 4400 -3195
rect 4800 -4795 5200 -3195
rect 5600 -4795 6000 -3195
rect 6400 -4795 6800 -3195
rect 7200 -4795 7600 -3195
rect 8000 -4795 8400 -3195
rect 8800 -4795 9200 -3195
rect 9600 -4795 10000 -3195
rect 10400 -4795 10800 -3195
rect 0 -7195 400 -5595
rect 800 -7195 1200 -5595
rect 1600 -7195 2000 -5595
rect 2400 -7195 2800 -5595
rect 3200 -7195 3600 -5595
rect 4000 -7195 4400 -5595
rect 4800 -7195 5200 -5595
rect 5600 -7195 6000 -5595
rect 6400 -7195 6800 -5595
rect 7200 -7195 7600 -5595
rect 8000 -7195 8400 -5595
rect 8800 -7195 9200 -5595
rect 9600 -7195 10000 -5595
rect 10400 -7195 10800 -5595
<< ndiff >>
rect -400 1585 0 1605
rect -400 25 -380 1585
rect -20 25 0 1585
rect -400 5 0 25
rect 400 1585 800 1605
rect 400 25 420 1585
rect 780 25 800 1585
rect 400 5 800 25
rect 1200 1585 1600 1605
rect 1200 25 1220 1585
rect 1580 25 1600 1585
rect 1200 5 1600 25
rect 2000 1585 2400 1605
rect 2000 25 2020 1585
rect 2380 25 2400 1585
rect 2000 5 2400 25
rect 2800 1585 3200 1605
rect 2800 25 2820 1585
rect 3180 25 3200 1585
rect 2800 5 3200 25
rect 3600 1585 4000 1605
rect 3600 25 3620 1585
rect 3980 25 4000 1585
rect 3600 5 4000 25
rect 4400 1585 4800 1605
rect 4400 25 4420 1585
rect 4780 25 4800 1585
rect 4400 5 4800 25
rect 5200 1585 5600 1605
rect 5200 25 5220 1585
rect 5580 25 5600 1585
rect 5200 5 5600 25
rect 6000 1585 6400 1605
rect 6000 25 6020 1585
rect 6380 25 6400 1585
rect 6000 5 6400 25
rect 6800 1585 7200 1605
rect 6800 25 6820 1585
rect 7180 25 7200 1585
rect 6800 5 7200 25
rect 7600 1585 8000 1605
rect 7600 25 7620 1585
rect 7980 25 8000 1585
rect 7600 5 8000 25
rect 8400 1585 8800 1605
rect 8400 25 8420 1585
rect 8780 25 8800 1585
rect 8400 5 8800 25
rect 9200 1585 9600 1605
rect 9200 25 9220 1585
rect 9580 25 9600 1585
rect 9200 5 9600 25
rect 10000 1585 10400 1605
rect 10000 25 10020 1585
rect 10380 25 10400 1585
rect 10000 5 10400 25
rect 10800 1585 11200 1605
rect 11600 1585 12000 1605
rect 10800 25 10820 1585
rect 11180 25 11200 1585
rect 11600 25 11620 1585
rect 11980 25 12000 1585
rect 10800 5 11200 25
rect 11600 5 12000 25
rect 12400 1585 12800 1605
rect 12400 25 12420 1585
rect 12780 25 12800 1585
rect 12400 5 12800 25
rect 13200 1585 13600 1605
rect 13200 25 13220 1585
rect 13580 25 13600 1585
rect 13200 5 13600 25
rect 14000 1585 14400 1605
rect 14000 25 14020 1585
rect 14380 25 14400 1585
rect 14000 5 14400 25
rect 14800 1585 15200 1605
rect 14800 25 14820 1585
rect 15180 25 15200 1585
rect 14800 5 15200 25
rect 15600 1585 16000 1605
rect 15600 25 15620 1585
rect 15980 25 16000 1585
rect 15600 5 16000 25
rect 16400 1585 16800 1605
rect 16400 25 16420 1585
rect 16780 25 16800 1585
rect 16400 5 16800 25
rect 17200 1585 17600 1605
rect 17200 25 17220 1585
rect 17580 25 17600 1585
rect 17200 5 17600 25
rect 18000 1585 18400 1605
rect 18000 25 18020 1585
rect 18380 25 18400 1585
rect 18000 5 18400 25
rect 18800 1585 19200 1605
rect 18800 25 18820 1585
rect 19180 25 19200 1585
rect 18800 5 19200 25
rect 19600 1585 20000 1605
rect 19600 25 19620 1585
rect 19980 25 20000 1585
rect 19600 5 20000 25
rect 20400 1585 20800 1605
rect 20400 25 20420 1585
rect 20780 25 20800 1585
rect 20400 5 20800 25
rect -400 -815 0 -795
rect -400 -2375 -380 -815
rect -20 -2375 0 -815
rect -400 -2395 0 -2375
rect 400 -815 800 -795
rect 400 -2375 420 -815
rect 780 -2375 800 -815
rect 400 -2395 800 -2375
rect 1200 -815 1600 -795
rect 1200 -2375 1220 -815
rect 1580 -2375 1600 -815
rect 1200 -2395 1600 -2375
rect 2000 -815 2400 -795
rect 2000 -2375 2020 -815
rect 2380 -2375 2400 -815
rect 2000 -2395 2400 -2375
rect 2800 -815 3200 -795
rect 2800 -2375 2820 -815
rect 3180 -2375 3200 -815
rect 2800 -2395 3200 -2375
rect 3600 -815 4000 -795
rect 3600 -2375 3620 -815
rect 3980 -2375 4000 -815
rect 3600 -2395 4000 -2375
rect 4400 -815 4800 -795
rect 4400 -2375 4420 -815
rect 4780 -2375 4800 -815
rect 4400 -2395 4800 -2375
rect 5200 -815 5600 -795
rect 5200 -2375 5220 -815
rect 5580 -2375 5600 -815
rect 5200 -2395 5600 -2375
rect 6000 -815 6400 -795
rect 6000 -2375 6020 -815
rect 6380 -2375 6400 -815
rect 6000 -2395 6400 -2375
rect 6800 -815 7200 -795
rect 6800 -2375 6820 -815
rect 7180 -2375 7200 -815
rect 6800 -2395 7200 -2375
rect 7600 -815 8000 -795
rect 7600 -2375 7620 -815
rect 7980 -2375 8000 -815
rect 7600 -2395 8000 -2375
rect 8400 -815 8800 -795
rect 8400 -2375 8420 -815
rect 8780 -2375 8800 -815
rect 8400 -2395 8800 -2375
rect 9200 -815 9600 -795
rect 9200 -2375 9220 -815
rect 9580 -2375 9600 -815
rect 9200 -2395 9600 -2375
rect 10000 -815 10400 -795
rect 10000 -2375 10020 -815
rect 10380 -2375 10400 -815
rect 10000 -2395 10400 -2375
rect 10800 -815 11200 -795
rect 10800 -2375 10820 -815
rect 11180 -2375 11200 -815
rect 10800 -2395 11200 -2375
rect -400 -3215 0 -3195
rect -400 -4775 -380 -3215
rect -20 -4775 0 -3215
rect -400 -4795 0 -4775
rect 400 -3215 800 -3195
rect 400 -4775 420 -3215
rect 780 -4775 800 -3215
rect 400 -4795 800 -4775
rect 1200 -3215 1600 -3195
rect 1200 -4775 1220 -3215
rect 1580 -4775 1600 -3215
rect 1200 -4795 1600 -4775
rect 2000 -3215 2400 -3195
rect 2000 -4775 2020 -3215
rect 2380 -4775 2400 -3215
rect 2000 -4795 2400 -4775
rect 2800 -3215 3200 -3195
rect 2800 -4775 2820 -3215
rect 3180 -4775 3200 -3215
rect 2800 -4795 3200 -4775
rect 3600 -3215 4000 -3195
rect 3600 -4775 3620 -3215
rect 3980 -4775 4000 -3215
rect 3600 -4795 4000 -4775
rect 4400 -3215 4800 -3195
rect 4400 -4775 4420 -3215
rect 4780 -4775 4800 -3215
rect 4400 -4795 4800 -4775
rect 5200 -3215 5600 -3195
rect 5200 -4775 5220 -3215
rect 5580 -4775 5600 -3215
rect 5200 -4795 5600 -4775
rect 6000 -3215 6400 -3195
rect 6000 -4775 6020 -3215
rect 6380 -4775 6400 -3215
rect 6000 -4795 6400 -4775
rect 6800 -3215 7200 -3195
rect 6800 -4775 6820 -3215
rect 7180 -4775 7200 -3215
rect 6800 -4795 7200 -4775
rect 7600 -3215 8000 -3195
rect 7600 -4775 7620 -3215
rect 7980 -4775 8000 -3215
rect 7600 -4795 8000 -4775
rect 8400 -3215 8800 -3195
rect 8400 -4775 8420 -3215
rect 8780 -4775 8800 -3215
rect 8400 -4795 8800 -4775
rect 9200 -3215 9600 -3195
rect 9200 -4775 9220 -3215
rect 9580 -4775 9600 -3215
rect 9200 -4795 9600 -4775
rect 10000 -3215 10400 -3195
rect 10000 -4775 10020 -3215
rect 10380 -4775 10400 -3215
rect 10000 -4795 10400 -4775
rect 10800 -3215 11200 -3195
rect 10800 -4775 10820 -3215
rect 11180 -4775 11200 -3215
rect 10800 -4795 11200 -4775
rect -400 -5615 0 -5595
rect -400 -7175 -380 -5615
rect -20 -7175 0 -5615
rect -400 -7195 0 -7175
rect 400 -5615 800 -5595
rect 400 -7175 420 -5615
rect 780 -7175 800 -5615
rect 400 -7195 800 -7175
rect 1200 -5615 1600 -5595
rect 1200 -7175 1220 -5615
rect 1580 -7175 1600 -5615
rect 1200 -7195 1600 -7175
rect 2000 -5615 2400 -5595
rect 2000 -7175 2020 -5615
rect 2380 -7175 2400 -5615
rect 2000 -7195 2400 -7175
rect 2800 -5615 3200 -5595
rect 2800 -7175 2820 -5615
rect 3180 -7175 3200 -5615
rect 2800 -7195 3200 -7175
rect 3600 -5615 4000 -5595
rect 3600 -7175 3620 -5615
rect 3980 -7175 4000 -5615
rect 3600 -7195 4000 -7175
rect 4400 -5615 4800 -5595
rect 4400 -7175 4420 -5615
rect 4780 -7175 4800 -5615
rect 4400 -7195 4800 -7175
rect 5200 -5615 5600 -5595
rect 5200 -7175 5220 -5615
rect 5580 -7175 5600 -5615
rect 5200 -7195 5600 -7175
rect 6000 -5615 6400 -5595
rect 6000 -7175 6020 -5615
rect 6380 -7175 6400 -5615
rect 6000 -7195 6400 -7175
rect 6800 -5615 7200 -5595
rect 6800 -7175 6820 -5615
rect 7180 -7175 7200 -5615
rect 6800 -7195 7200 -7175
rect 7600 -5615 8000 -5595
rect 7600 -7175 7620 -5615
rect 7980 -7175 8000 -5615
rect 7600 -7195 8000 -7175
rect 8400 -5615 8800 -5595
rect 8400 -7175 8420 -5615
rect 8780 -7175 8800 -5615
rect 8400 -7195 8800 -7175
rect 9200 -5615 9600 -5595
rect 9200 -7175 9220 -5615
rect 9580 -7175 9600 -5615
rect 9200 -7195 9600 -7175
rect 10000 -5615 10400 -5595
rect 10000 -7175 10020 -5615
rect 10380 -7175 10400 -5615
rect 10000 -7195 10400 -7175
rect 10800 -5615 11200 -5595
rect 10800 -7175 10820 -5615
rect 11180 -7175 11200 -5615
rect 10800 -7195 11200 -7175
<< ndiffc >>
rect -380 25 -20 1585
rect 420 25 780 1585
rect 1220 25 1580 1585
rect 2020 25 2380 1585
rect 2820 25 3180 1585
rect 3620 25 3980 1585
rect 4420 25 4780 1585
rect 5220 25 5580 1585
rect 6020 25 6380 1585
rect 6820 25 7180 1585
rect 7620 25 7980 1585
rect 8420 25 8780 1585
rect 9220 25 9580 1585
rect 10020 25 10380 1585
rect 10820 25 11180 1585
rect 11620 25 11980 1585
rect 12420 25 12780 1585
rect 13220 25 13580 1585
rect 14020 25 14380 1585
rect 14820 25 15180 1585
rect 15620 25 15980 1585
rect 16420 25 16780 1585
rect 17220 25 17580 1585
rect 18020 25 18380 1585
rect 18820 25 19180 1585
rect 19620 25 19980 1585
rect 20420 25 20780 1585
rect -380 -2375 -20 -815
rect 420 -2375 780 -815
rect 1220 -2375 1580 -815
rect 2020 -2375 2380 -815
rect 2820 -2375 3180 -815
rect 3620 -2375 3980 -815
rect 4420 -2375 4780 -815
rect 5220 -2375 5580 -815
rect 6020 -2375 6380 -815
rect 6820 -2375 7180 -815
rect 7620 -2375 7980 -815
rect 8420 -2375 8780 -815
rect 9220 -2375 9580 -815
rect 10020 -2375 10380 -815
rect 10820 -2375 11180 -815
rect -380 -4775 -20 -3215
rect 420 -4775 780 -3215
rect 1220 -4775 1580 -3215
rect 2020 -4775 2380 -3215
rect 2820 -4775 3180 -3215
rect 3620 -4775 3980 -3215
rect 4420 -4775 4780 -3215
rect 5220 -4775 5580 -3215
rect 6020 -4775 6380 -3215
rect 6820 -4775 7180 -3215
rect 7620 -4775 7980 -3215
rect 8420 -4775 8780 -3215
rect 9220 -4775 9580 -3215
rect 10020 -4775 10380 -3215
rect 10820 -4775 11180 -3215
rect -380 -7175 -20 -5615
rect 420 -7175 780 -5615
rect 1220 -7175 1580 -5615
rect 2020 -7175 2380 -5615
rect 2820 -7175 3180 -5615
rect 3620 -7175 3980 -5615
rect 4420 -7175 4780 -5615
rect 5220 -7175 5580 -5615
rect 6020 -7175 6380 -5615
rect 6820 -7175 7180 -5615
rect 7620 -7175 7980 -5615
rect 8420 -7175 8780 -5615
rect 9220 -7175 9580 -5615
rect 10020 -7175 10380 -5615
rect 10820 -7175 11180 -5615
<< psubdiff >>
rect -800 1585 -400 1605
rect -800 25 -780 1585
rect -420 25 -400 1585
rect -800 5 -400 25
rect 11200 1585 11600 1605
rect 11200 25 11220 1585
rect 11580 25 11600 1585
rect 11200 5 11600 25
rect 20800 1585 21200 1605
rect 20800 25 20820 1585
rect 21180 25 21200 1585
rect 20800 5 21200 25
rect -800 -815 -400 -795
rect -800 -2375 -780 -815
rect -420 -2375 -400 -815
rect -800 -2395 -400 -2375
rect -800 -3215 -400 -3195
rect -800 -4775 -780 -3215
rect -420 -4775 -400 -3215
rect -800 -4795 -400 -4775
rect -800 -5615 -400 -5595
rect -800 -7175 -780 -5615
rect -420 -7175 -400 -5615
rect -800 -7195 -400 -7175
<< psubdiffcont >>
rect -780 25 -420 1585
rect 11220 25 11580 1585
rect 20820 25 21180 1585
rect -780 -2375 -420 -815
rect -780 -4775 -420 -3215
rect -780 -7175 -420 -5615
<< poly >>
rect 0 1605 400 1620
rect 800 1605 1200 1620
rect 1600 1605 2000 1620
rect 2400 1605 2800 1620
rect 3200 1605 3600 1620
rect 4000 1605 4400 1620
rect 4800 1605 5200 1620
rect 5600 1605 6000 1620
rect 6400 1605 6800 1620
rect 7200 1605 7600 1620
rect 8000 1605 8400 1620
rect 8800 1605 9200 1620
rect 9600 1605 10000 1620
rect 10400 1605 10800 1620
rect 12000 1605 12400 1620
rect 12800 1605 13200 1620
rect 13600 1605 14000 1620
rect 14400 1605 14800 1620
rect 15200 1605 15600 1620
rect 16000 1605 16400 1620
rect 16800 1605 17200 1620
rect 17600 1605 18000 1620
rect 18400 1605 18800 1620
rect 19200 1605 19600 1620
rect 20000 1605 20400 1620
rect 0 -10 400 5
rect 800 -10 1200 5
rect 1600 -10 2000 5
rect 2400 -10 2800 5
rect 3200 -10 3600 5
rect 4000 -10 4400 5
rect 4800 -10 5200 5
rect 5600 -10 6000 5
rect 6400 -10 6800 5
rect 7200 -10 7600 5
rect 8000 -10 8400 5
rect 8800 -10 9200 5
rect 9600 -10 10000 5
rect 10400 -10 10800 5
rect 12000 -10 12400 5
rect 12800 -10 13200 5
rect 13600 -10 14000 5
rect 14400 -10 14800 5
rect 15200 -10 15600 5
rect 16000 -10 16400 5
rect 16800 -10 17200 5
rect 17600 -10 18000 5
rect 18400 -10 18800 5
rect 19200 -10 19600 5
rect 20000 -10 20400 5
rect -390 -20 1200 -10
rect -390 -100 -380 -20
rect -20 -100 420 -20
rect 780 -100 1200 -20
rect -390 -110 1200 -100
rect 9600 -20 11190 -10
rect 9600 -100 10020 -20
rect 10380 -100 10820 -20
rect 11180 -100 11190 -20
rect 9600 -110 11190 -100
rect 11610 -20 12400 -10
rect 11610 -100 11620 -20
rect 11980 -100 12400 -20
rect 11610 -110 12400 -100
rect 20000 -20 20790 -10
rect 20000 -100 20420 -20
rect 20780 -100 20790 -20
rect 20000 -110 20790 -100
rect 0 -795 400 -780
rect 800 -795 1200 -780
rect 1600 -795 2000 -780
rect 2400 -795 2800 -780
rect 3200 -795 3600 -780
rect 4000 -795 4400 -780
rect 4800 -795 5200 -780
rect 5600 -795 6000 -780
rect 6400 -795 6800 -780
rect 7200 -795 7600 -780
rect 8000 -795 8400 -780
rect 8800 -795 9200 -780
rect 9600 -795 10000 -780
rect 10400 -795 10800 -780
rect 0 -2410 400 -2395
rect 800 -2410 1200 -2395
rect 1600 -2410 2000 -2395
rect 2400 -2410 2800 -2395
rect 3200 -2410 3600 -2395
rect 4000 -2410 4400 -2395
rect 4800 -2410 5200 -2395
rect 5600 -2410 6000 -2395
rect 6400 -2410 6800 -2395
rect 7200 -2410 7600 -2395
rect 8000 -2410 8400 -2395
rect 8800 -2410 9200 -2395
rect 9600 -2410 10000 -2395
rect 10400 -2410 10800 -2395
rect -390 -2420 1200 -2410
rect -390 -2500 -380 -2420
rect -20 -2500 420 -2420
rect 780 -2500 1200 -2420
rect -390 -2510 1200 -2500
rect 9600 -2420 11190 -2410
rect 9600 -2500 10020 -2420
rect 10380 -2500 10820 -2420
rect 11180 -2500 11190 -2420
rect 9600 -2510 11190 -2500
rect 0 -3195 400 -3180
rect 800 -3195 1200 -3180
rect 1600 -3195 2000 -3180
rect 2400 -3195 2800 -3180
rect 3200 -3195 3600 -3180
rect 4000 -3195 4400 -3180
rect 4800 -3195 5200 -3180
rect 5600 -3195 6000 -3180
rect 6400 -3195 6800 -3180
rect 7200 -3195 7600 -3180
rect 8000 -3195 8400 -3180
rect 8800 -3195 9200 -3180
rect 9600 -3195 10000 -3180
rect 10400 -3195 10800 -3180
rect 0 -4810 400 -4795
rect 800 -4810 1200 -4795
rect 1600 -4810 2000 -4795
rect 2400 -4810 2800 -4795
rect 3200 -4810 3600 -4795
rect 4000 -4810 4400 -4795
rect 4800 -4810 5200 -4795
rect 5600 -4810 6000 -4795
rect 6400 -4810 6800 -4795
rect 7200 -4810 7600 -4795
rect 8000 -4810 8400 -4795
rect 8800 -4810 9200 -4795
rect 9600 -4810 10000 -4795
rect 10400 -4810 10800 -4795
rect -390 -4820 400 -4810
rect -390 -4900 -380 -4820
rect -20 -4900 400 -4820
rect -390 -4910 400 -4900
rect 10400 -4820 11190 -4810
rect 10400 -4900 10820 -4820
rect 11180 -4900 11190 -4820
rect 10400 -4910 11190 -4900
rect 0 -5595 400 -5580
rect 800 -5595 1200 -5580
rect 1600 -5595 2000 -5580
rect 2400 -5595 2800 -5580
rect 3200 -5595 3600 -5580
rect 4000 -5595 4400 -5580
rect 4800 -5595 5200 -5580
rect 5600 -5595 6000 -5580
rect 6400 -5595 6800 -5580
rect 7200 -5595 7600 -5580
rect 8000 -5595 8400 -5580
rect 8800 -5595 9200 -5580
rect 9600 -5595 10000 -5580
rect 10400 -5595 10800 -5580
rect 0 -7210 400 -7195
rect 800 -7210 1200 -7195
rect 1600 -7210 2000 -7195
rect 2400 -7210 2800 -7195
rect 3200 -7210 3600 -7195
rect 4000 -7210 4400 -7195
rect 4800 -7210 5200 -7195
rect 5600 -7210 6000 -7195
rect 6400 -7210 6800 -7195
rect 7200 -7210 7600 -7195
rect 8000 -7210 8400 -7195
rect 8800 -7210 9200 -7195
rect 9600 -7210 10000 -7195
rect 10400 -7210 10800 -7195
rect -390 -7220 400 -7210
rect -390 -7300 -380 -7220
rect -20 -7300 400 -7220
rect -390 -7310 400 -7300
rect 10400 -7220 11190 -7210
rect 10400 -7300 10820 -7220
rect 11180 -7300 11190 -7220
rect 10400 -7310 11190 -7300
<< polycont >>
rect -380 -100 -20 -20
rect 420 -100 780 -20
rect 10020 -100 10380 -20
rect 10820 -100 11180 -20
rect 11620 -100 11980 -20
rect 20420 -100 20780 -20
rect -380 -2500 -20 -2420
rect 420 -2500 780 -2420
rect 10020 -2500 10380 -2420
rect 10820 -2500 11180 -2420
rect -380 -4900 -20 -4820
rect 10820 -4900 11180 -4820
rect -380 -7300 -20 -7220
rect 10820 -7300 11180 -7220
<< locali >>
rect -790 1585 -10 1595
rect -790 25 -780 1585
rect -420 25 -380 1585
rect -20 25 -10 1585
rect -790 15 -10 25
rect -390 -20 -10 15
rect -390 -100 -380 -20
rect -20 -100 -10 -20
rect -390 -110 -10 -100
rect 410 1585 790 1595
rect 410 25 420 1585
rect 780 25 790 1585
rect 410 -20 790 25
rect 1210 1585 1590 1595
rect 1210 25 1220 1585
rect 1580 25 1590 1585
rect 1210 15 1590 25
rect 2010 1585 2390 1595
rect 2010 25 2020 1585
rect 2380 25 2390 1585
rect 2010 15 2390 25
rect 2810 1585 3190 1595
rect 2810 25 2820 1585
rect 3180 25 3190 1585
rect 2810 15 3190 25
rect 3610 1585 3990 1595
rect 3610 25 3620 1585
rect 3980 25 3990 1585
rect 3610 15 3990 25
rect 4410 1585 4790 1595
rect 4410 25 4420 1585
rect 4780 25 4790 1585
rect 4410 15 4790 25
rect 5210 1585 5590 1595
rect 5210 25 5220 1585
rect 5580 25 5590 1585
rect 5210 15 5590 25
rect 6010 1585 6390 1595
rect 6010 25 6020 1585
rect 6380 25 6390 1585
rect 6010 15 6390 25
rect 6810 1585 7190 1595
rect 6810 25 6820 1585
rect 7180 25 7190 1585
rect 6810 15 7190 25
rect 7610 1585 7990 1595
rect 7610 25 7620 1585
rect 7980 25 7990 1585
rect 7610 15 7990 25
rect 8410 1585 8790 1595
rect 8410 25 8420 1585
rect 8780 25 8790 1585
rect 8410 15 8790 25
rect 9210 1585 9590 1595
rect 9210 25 9220 1585
rect 9580 25 9590 1585
rect 9210 15 9590 25
rect 10010 1585 10390 1595
rect 10010 25 10020 1585
rect 10380 25 10390 1585
rect 410 -100 420 -20
rect 780 -100 790 -20
rect 410 -110 790 -100
rect 10010 -20 10390 25
rect 10010 -100 10020 -20
rect 10380 -100 10390 -20
rect 10010 -110 10390 -100
rect 10810 1585 11990 1595
rect 10810 25 10820 1585
rect 11180 25 11220 1585
rect 11580 25 11620 1585
rect 11980 25 11990 1585
rect 10810 15 11990 25
rect 12410 1585 12790 1595
rect 12410 25 12420 1585
rect 12780 25 12790 1585
rect 12410 15 12790 25
rect 13210 1585 13590 1595
rect 13210 25 13220 1585
rect 13580 25 13590 1585
rect 13210 15 13590 25
rect 14010 1585 14390 1595
rect 14010 25 14020 1585
rect 14380 25 14390 1585
rect 14010 15 14390 25
rect 14810 1585 15190 1595
rect 14810 25 14820 1585
rect 15180 25 15190 1585
rect 14810 15 15190 25
rect 15610 1585 15990 1595
rect 15610 25 15620 1585
rect 15980 25 15990 1585
rect 15610 15 15990 25
rect 16410 1585 16790 1595
rect 16410 25 16420 1585
rect 16780 25 16790 1585
rect 16410 15 16790 25
rect 17210 1585 17590 1595
rect 17210 25 17220 1585
rect 17580 25 17590 1585
rect 17210 15 17590 25
rect 18010 1585 18390 1595
rect 18010 25 18020 1585
rect 18380 25 18390 1585
rect 18010 15 18390 25
rect 18810 1585 19190 1595
rect 18810 25 18820 1585
rect 19180 25 19190 1585
rect 18810 15 19190 25
rect 19610 1585 19990 1595
rect 19610 25 19620 1585
rect 19980 25 19990 1585
rect 19610 15 19990 25
rect 20410 1585 21190 1595
rect 20410 25 20420 1585
rect 20780 25 20820 1585
rect 21180 25 21190 1585
rect 20410 15 21190 25
rect 10810 -20 11190 15
rect 10810 -100 10820 -20
rect 11180 -100 11190 -20
rect 10810 -110 11190 -100
rect 11610 -20 11990 15
rect 11610 -100 11620 -20
rect 11980 -100 11990 -20
rect 11610 -110 11990 -100
rect 20410 -20 20790 15
rect 20410 -100 20420 -20
rect 20780 -100 20790 -20
rect 20410 -110 20790 -100
rect -790 -815 -10 -805
rect -790 -2375 -780 -815
rect -420 -2375 -380 -815
rect -20 -2375 -10 -815
rect -790 -2385 -10 -2375
rect -390 -2420 -10 -2385
rect -390 -2500 -380 -2420
rect -20 -2500 -10 -2420
rect -390 -2510 -10 -2500
rect 410 -815 790 -805
rect 410 -2375 420 -815
rect 780 -2375 790 -815
rect 410 -2420 790 -2375
rect 1210 -815 1590 -805
rect 1210 -2375 1220 -815
rect 1580 -2375 1590 -815
rect 1210 -2385 1590 -2375
rect 2010 -815 2390 -805
rect 2010 -2375 2020 -815
rect 2380 -2375 2390 -815
rect 2010 -2385 2390 -2375
rect 2810 -815 3190 -805
rect 2810 -2375 2820 -815
rect 3180 -2375 3190 -815
rect 2810 -2385 3190 -2375
rect 3610 -815 3990 -805
rect 3610 -2375 3620 -815
rect 3980 -2375 3990 -815
rect 3610 -2385 3990 -2375
rect 4410 -815 4790 -805
rect 4410 -2375 4420 -815
rect 4780 -2375 4790 -815
rect 4410 -2385 4790 -2375
rect 5210 -815 5590 -805
rect 5210 -2375 5220 -815
rect 5580 -2375 5590 -815
rect 5210 -2385 5590 -2375
rect 6010 -815 6390 -805
rect 6010 -2375 6020 -815
rect 6380 -2375 6390 -815
rect 6010 -2385 6390 -2375
rect 6810 -815 7190 -805
rect 6810 -2375 6820 -815
rect 7180 -2375 7190 -815
rect 6810 -2385 7190 -2375
rect 7610 -815 7990 -805
rect 7610 -2375 7620 -815
rect 7980 -2375 7990 -815
rect 7610 -2385 7990 -2375
rect 8410 -815 8790 -805
rect 8410 -2375 8420 -815
rect 8780 -2375 8790 -815
rect 8410 -2385 8790 -2375
rect 9210 -815 9590 -805
rect 9210 -2375 9220 -815
rect 9580 -2375 9590 -815
rect 9210 -2385 9590 -2375
rect 10010 -815 10390 -805
rect 10010 -2375 10020 -815
rect 10380 -2375 10390 -815
rect 410 -2500 420 -2420
rect 780 -2500 790 -2420
rect 410 -2510 790 -2500
rect 10010 -2420 10390 -2375
rect 10010 -2500 10020 -2420
rect 10380 -2500 10390 -2420
rect 10010 -2510 10390 -2500
rect 10810 -815 11200 -805
rect 10810 -2375 10820 -815
rect 11180 -2375 11200 -815
rect 10810 -2385 11200 -2375
rect 10810 -2420 11190 -2385
rect 10810 -2500 10820 -2420
rect 11180 -2500 11190 -2420
rect 10810 -2510 11190 -2500
rect -790 -3215 -10 -3205
rect -790 -4775 -780 -3215
rect -420 -4775 -380 -3215
rect -20 -4775 -10 -3215
rect -790 -4785 -10 -4775
rect 410 -3215 790 -3205
rect 410 -4775 420 -3215
rect 780 -4775 790 -3215
rect 410 -4785 790 -4775
rect 1210 -3215 1590 -3205
rect 1210 -4775 1220 -3215
rect 1580 -4775 1590 -3215
rect 1210 -4785 1590 -4775
rect 2010 -3215 2390 -3205
rect 2010 -4775 2020 -3215
rect 2380 -4775 2390 -3215
rect 2010 -4785 2390 -4775
rect 2810 -3215 3190 -3205
rect 2810 -4775 2820 -3215
rect 3180 -4775 3190 -3215
rect 2810 -4785 3190 -4775
rect 3610 -3215 3990 -3205
rect 3610 -4775 3620 -3215
rect 3980 -4775 3990 -3215
rect 3610 -4785 3990 -4775
rect 4410 -3215 4790 -3205
rect 4410 -4775 4420 -3215
rect 4780 -4775 4790 -3215
rect 4410 -4785 4790 -4775
rect 5210 -3215 5590 -3205
rect 5210 -4775 5220 -3215
rect 5580 -4775 5590 -3215
rect 5210 -4785 5590 -4775
rect 6010 -3215 6390 -3205
rect 6010 -4775 6020 -3215
rect 6380 -4775 6390 -3215
rect 6010 -4785 6390 -4775
rect 6810 -3215 7190 -3205
rect 6810 -4775 6820 -3215
rect 7180 -4775 7190 -3215
rect 6810 -4785 7190 -4775
rect 7610 -3215 7990 -3205
rect 7610 -4775 7620 -3215
rect 7980 -4775 7990 -3215
rect 7610 -4785 7990 -4775
rect 8410 -3215 8790 -3205
rect 8410 -4775 8420 -3215
rect 8780 -4775 8790 -3215
rect 8410 -4785 8790 -4775
rect 9210 -3215 9590 -3205
rect 9210 -4775 9220 -3215
rect 9580 -4775 9590 -3215
rect 9210 -4785 9590 -4775
rect 10010 -3215 10390 -3205
rect 10010 -4775 10020 -3215
rect 10380 -4775 10390 -3215
rect 10010 -4785 10390 -4775
rect 10810 -3215 11200 -3205
rect 10810 -4775 10820 -3215
rect 11180 -4775 11200 -3215
rect 10810 -4785 11200 -4775
rect -390 -4820 -10 -4785
rect -390 -4900 -380 -4820
rect -20 -4900 -10 -4820
rect -390 -4910 -10 -4900
rect 10810 -4820 11190 -4785
rect 10810 -4900 10820 -4820
rect 11180 -4900 11190 -4820
rect 10810 -4910 11190 -4900
rect -790 -5615 -10 -5605
rect -790 -7175 -780 -5615
rect -420 -7175 -380 -5615
rect -20 -7175 -10 -5615
rect -790 -7185 -10 -7175
rect 410 -5615 790 -5605
rect 410 -7175 420 -5615
rect 780 -7175 790 -5615
rect 410 -7185 790 -7175
rect 1210 -5615 1590 -5605
rect 1210 -7175 1220 -5615
rect 1580 -7175 1590 -5615
rect 1210 -7185 1590 -7175
rect 2010 -5615 2390 -5605
rect 2010 -7175 2020 -5615
rect 2380 -7175 2390 -5615
rect 2010 -7185 2390 -7175
rect 2810 -5615 3190 -5605
rect 2810 -7175 2820 -5615
rect 3180 -7175 3190 -5615
rect 2810 -7185 3190 -7175
rect 3610 -5615 3990 -5605
rect 3610 -7175 3620 -5615
rect 3980 -7175 3990 -5615
rect 3610 -7185 3990 -7175
rect 4410 -5615 4790 -5605
rect 4410 -7175 4420 -5615
rect 4780 -7175 4790 -5615
rect 4410 -7185 4790 -7175
rect 5210 -5615 5590 -5605
rect 5210 -7175 5220 -5615
rect 5580 -7175 5590 -5615
rect 5210 -7185 5590 -7175
rect 6010 -5615 6390 -5605
rect 6010 -7175 6020 -5615
rect 6380 -7175 6390 -5615
rect 6010 -7185 6390 -7175
rect 6810 -5615 7190 -5605
rect 6810 -7175 6820 -5615
rect 7180 -7175 7190 -5615
rect 6810 -7185 7190 -7175
rect 7610 -5615 7990 -5605
rect 7610 -7175 7620 -5615
rect 7980 -7175 7990 -5615
rect 7610 -7185 7990 -7175
rect 8410 -5615 8790 -5605
rect 8410 -7175 8420 -5615
rect 8780 -7175 8790 -5615
rect 8410 -7185 8790 -7175
rect 9210 -5615 9590 -5605
rect 9210 -7175 9220 -5615
rect 9580 -7175 9590 -5615
rect 9210 -7185 9590 -7175
rect 10010 -5615 10390 -5605
rect 10010 -7175 10020 -5615
rect 10380 -7175 10390 -5615
rect 10010 -7185 10390 -7175
rect 10810 -5615 11200 -5605
rect 10810 -7175 10820 -5615
rect 11180 -7175 11200 -5615
rect 10810 -7185 11200 -7175
rect -390 -7220 -10 -7185
rect -390 -7300 -380 -7220
rect -20 -7300 -10 -7220
rect -390 -7310 -10 -7300
rect 10810 -7220 11190 -7185
rect 10810 -7300 10820 -7220
rect 11180 -7300 11190 -7220
rect 10810 -7310 11190 -7300
<< end >>
